magic
tech scmos
timestamp 1764608577
<< nwell >>
rect 26 342 74 363
rect 17 285 74 342
rect 32 261 74 285
rect 194 270 231 301
rect 167 267 231 270
rect -1 226 36 253
rect -2 223 36 226
rect 167 223 232 267
rect 323 245 371 266
rect -2 187 35 223
rect 314 188 371 245
rect 329 164 371 188
rect 23 135 71 156
rect 14 78 71 135
rect 29 54 71 78
rect 2 13 45 48
rect 2 -20 42 13
<< ntransistor >>
rect 82 345 92 347
rect 80 329 100 331
rect 80 321 100 323
rect 80 313 100 315
rect 80 304 100 306
rect 237 283 247 285
rect 82 280 92 282
rect 240 254 260 256
rect 379 248 389 250
rect 240 244 260 246
rect 42 235 52 237
rect 240 234 260 236
rect 377 232 397 234
rect 377 224 397 226
rect 377 216 397 218
rect 41 210 51 212
rect 377 207 397 209
rect 41 198 51 200
rect 379 183 389 185
rect 79 138 89 140
rect 77 122 97 124
rect 77 114 97 116
rect 77 106 97 108
rect 77 97 97 99
rect 79 73 89 75
rect 51 27 61 29
rect 49 -1 69 1
rect 49 -9 69 -7
<< ptransistor >>
rect 43 345 63 347
rect 23 329 63 331
rect 23 321 63 323
rect 23 313 63 315
rect 23 304 63 306
rect 205 283 225 285
rect 43 280 63 282
rect 186 254 226 256
rect 340 248 360 250
rect 186 244 226 246
rect 10 235 30 237
rect 186 234 226 236
rect 320 232 360 234
rect 320 224 360 226
rect 320 216 360 218
rect 9 210 29 212
rect 320 207 360 209
rect 9 198 29 200
rect 340 183 360 185
rect 40 138 60 140
rect 20 122 60 124
rect 20 114 60 116
rect 20 106 60 108
rect 20 97 60 99
rect 40 73 60 75
rect 19 27 39 29
rect 16 -1 36 1
rect 16 -9 36 -7
<< ndiffusion >>
rect 82 349 84 353
rect 88 349 92 353
rect 82 347 92 349
rect 82 344 92 345
rect 82 340 88 344
rect 84 332 100 336
rect 80 331 100 332
rect 80 323 100 329
rect 80 320 100 321
rect 80 316 96 320
rect 80 315 100 316
rect 80 306 100 313
rect 80 303 100 304
rect 84 299 100 303
rect 86 283 92 287
rect 237 286 239 290
rect 243 286 247 290
rect 237 285 247 286
rect 82 282 92 283
rect 82 278 92 280
rect 237 282 247 283
rect 237 278 243 282
rect 82 274 88 278
rect 240 257 256 261
rect 240 256 260 257
rect 240 252 260 254
rect 244 248 260 252
rect 240 246 260 248
rect 379 252 381 256
rect 385 252 389 256
rect 379 250 389 252
rect 42 238 44 242
rect 48 238 52 242
rect 42 237 52 238
rect 42 234 52 235
rect 42 230 48 234
rect 240 236 260 244
rect 379 247 389 248
rect 379 243 385 247
rect 240 233 260 234
rect 240 229 256 233
rect 381 235 397 239
rect 377 234 397 235
rect 377 226 397 232
rect 45 213 51 217
rect 377 223 397 224
rect 377 219 393 223
rect 377 218 397 219
rect 41 212 51 213
rect 41 200 51 210
rect 377 209 397 216
rect 377 206 397 207
rect 381 202 397 206
rect 41 197 51 198
rect 41 193 47 197
rect 383 186 389 190
rect 379 185 389 186
rect 379 181 389 183
rect 379 177 385 181
rect 79 142 81 146
rect 85 142 89 146
rect 79 140 89 142
rect 79 137 89 138
rect 79 133 85 137
rect 81 125 97 129
rect 77 124 97 125
rect 77 116 97 122
rect 77 113 97 114
rect 77 109 93 113
rect 77 108 97 109
rect 77 99 97 106
rect 77 96 97 97
rect 81 92 97 96
rect 83 76 89 80
rect 79 75 89 76
rect 79 71 89 73
rect 79 67 85 71
rect 51 30 53 34
rect 57 30 61 34
rect 51 29 61 30
rect 51 26 61 27
rect 51 22 57 26
rect 49 1 69 2
rect 49 -2 69 -1
rect 49 -7 69 -6
rect 49 -10 69 -9
<< pdiffusion >>
rect 43 349 57 353
rect 61 349 63 353
rect 43 347 63 349
rect 43 344 63 345
rect 43 340 59 344
rect 43 339 63 340
rect 27 332 63 336
rect 23 331 63 332
rect 23 328 63 329
rect 23 324 59 328
rect 23 323 63 324
rect 23 320 63 321
rect 27 316 63 320
rect 23 315 63 316
rect 23 311 63 313
rect 23 307 59 311
rect 23 306 63 307
rect 23 303 63 304
rect 27 299 63 303
rect 43 287 63 288
rect 43 283 59 287
rect 43 282 63 283
rect 205 286 219 290
rect 223 286 225 290
rect 205 285 225 286
rect 205 282 225 283
rect 43 278 63 280
rect 43 274 59 278
rect 209 278 225 282
rect 186 257 222 261
rect 186 256 226 257
rect 186 252 226 254
rect 186 248 222 252
rect 186 246 226 248
rect 340 252 354 256
rect 358 252 360 256
rect 340 250 360 252
rect 340 247 360 248
rect 186 242 226 244
rect 10 238 24 242
rect 28 238 30 242
rect 10 237 30 238
rect 190 238 226 242
rect 10 234 30 235
rect 14 230 30 234
rect 186 236 226 238
rect 340 243 356 247
rect 340 242 360 243
rect 324 235 360 239
rect 186 233 226 234
rect 186 229 222 233
rect 320 234 360 235
rect 320 231 360 232
rect 320 227 356 231
rect 320 226 360 227
rect 320 223 360 224
rect 324 219 360 223
rect 13 213 29 217
rect 9 212 29 213
rect 320 218 360 219
rect 320 214 360 216
rect 320 210 356 214
rect 9 207 29 210
rect 9 203 24 207
rect 28 203 29 207
rect 9 200 29 203
rect 320 209 360 210
rect 320 206 360 207
rect 324 202 360 206
rect 9 197 29 198
rect 13 193 29 197
rect 340 190 360 191
rect 340 186 356 190
rect 340 185 360 186
rect 340 181 360 183
rect 340 177 356 181
rect 40 142 54 146
rect 58 142 60 146
rect 40 140 60 142
rect 40 137 60 138
rect 40 133 56 137
rect 40 132 60 133
rect 24 125 60 129
rect 20 124 60 125
rect 20 121 60 122
rect 20 117 56 121
rect 20 116 60 117
rect 20 113 60 114
rect 24 109 60 113
rect 20 108 60 109
rect 20 104 60 106
rect 20 100 56 104
rect 20 99 60 100
rect 20 96 60 97
rect 24 92 60 96
rect 40 80 60 81
rect 40 76 56 80
rect 40 75 60 76
rect 40 71 60 73
rect 40 67 56 71
rect 19 30 33 34
rect 37 30 39 34
rect 19 29 39 30
rect 19 26 39 27
rect 23 22 39 26
rect 16 1 36 2
rect 16 -2 36 -1
rect 16 -7 36 -6
rect 16 -10 36 -9
<< ndcontact >>
rect 84 349 88 353
rect 88 340 92 344
rect 80 332 84 336
rect 96 316 100 320
rect 80 299 84 303
rect 82 283 86 287
rect 239 286 243 290
rect 243 278 247 282
rect 88 274 92 278
rect 256 257 260 261
rect 240 248 244 252
rect 381 252 385 256
rect 44 238 48 242
rect 48 230 52 234
rect 385 243 389 247
rect 256 229 260 233
rect 377 235 381 239
rect 41 213 45 217
rect 393 219 397 223
rect 377 202 381 206
rect 47 193 51 197
rect 379 186 383 190
rect 385 177 389 181
rect 81 142 85 146
rect 85 133 89 137
rect 77 125 81 129
rect 93 109 97 113
rect 77 92 81 96
rect 79 76 83 80
rect 85 67 89 71
rect 53 30 57 34
rect 57 22 61 26
rect 49 2 69 6
rect 49 -6 69 -2
rect 49 -14 69 -10
<< pdcontact >>
rect 57 349 61 353
rect 59 340 63 344
rect 23 332 27 336
rect 59 324 63 328
rect 23 316 27 320
rect 117 316 121 320
rect 59 307 63 311
rect 23 299 27 303
rect 59 283 63 287
rect 219 286 223 290
rect 59 274 63 278
rect 205 278 209 282
rect 222 257 226 261
rect 222 248 226 252
rect 354 252 358 256
rect 24 238 28 242
rect 186 238 190 242
rect 10 230 14 234
rect 356 243 360 247
rect 320 235 324 239
rect 222 229 226 233
rect 356 227 360 231
rect 320 219 324 223
rect 9 213 13 217
rect 414 219 418 223
rect 356 210 360 214
rect 24 203 28 207
rect 320 202 324 206
rect 9 193 13 197
rect 356 186 360 190
rect 356 177 360 181
rect 54 142 58 146
rect 56 133 60 137
rect 20 125 24 129
rect 56 117 60 121
rect 20 109 24 113
rect 114 109 118 113
rect 56 100 60 104
rect 20 92 24 96
rect 56 76 60 80
rect 56 67 60 71
rect 33 30 37 34
rect 19 22 23 26
rect 16 2 36 6
rect 16 -6 36 -2
rect 16 -14 36 -10
<< psubstratepcontact >>
rect 104 316 108 320
rect 251 278 255 282
rect 56 230 60 234
rect 264 238 268 242
rect 401 219 405 223
rect 55 193 59 197
rect 101 109 105 113
rect 65 22 69 26
rect 73 -14 77 -10
<< nsubstratencontact >>
rect 197 278 201 282
rect 59 264 63 268
rect 178 238 182 242
rect 2 230 6 234
rect 1 203 5 207
rect 356 167 360 171
rect 56 57 60 61
rect 11 22 15 26
rect 7 -14 11 -10
<< polysilicon >>
rect 42 345 43 347
rect 63 345 82 347
rect 92 345 95 347
rect -5 329 23 331
rect 63 329 80 331
rect 100 329 103 331
rect 11 321 23 323
rect 63 321 80 323
rect 100 321 103 323
rect -6 313 23 315
rect 63 313 80 315
rect 100 313 103 315
rect -5 304 23 306
rect 63 304 80 306
rect 100 304 103 306
rect 202 283 205 285
rect 225 283 237 285
rect 247 283 250 285
rect 42 280 43 282
rect 63 280 82 282
rect 92 280 95 282
rect 175 254 186 256
rect 226 254 240 256
rect 260 254 263 256
rect 339 248 340 250
rect 360 248 379 250
rect 389 248 392 250
rect 175 244 186 246
rect 226 244 240 246
rect 260 244 263 246
rect 7 235 10 237
rect 30 235 42 237
rect 52 235 55 237
rect 175 234 186 236
rect 226 234 240 236
rect 260 234 263 236
rect 292 232 320 234
rect 360 232 377 234
rect 397 232 400 234
rect 308 224 320 226
rect 360 224 377 226
rect 397 224 400 226
rect 291 216 320 218
rect 360 216 377 218
rect 397 216 400 218
rect -2 210 9 212
rect 29 210 41 212
rect 51 210 54 212
rect 292 207 320 209
rect 360 207 377 209
rect 397 207 400 209
rect -2 198 9 200
rect 29 198 41 200
rect 51 198 54 200
rect 339 183 340 185
rect 360 183 379 185
rect 389 183 392 185
rect 39 138 40 140
rect 60 138 79 140
rect 89 138 92 140
rect -8 122 20 124
rect 60 122 77 124
rect 97 122 100 124
rect 8 114 20 116
rect 60 114 77 116
rect 97 114 100 116
rect -9 106 20 108
rect 60 106 77 108
rect 97 106 100 108
rect -8 97 20 99
rect 60 97 77 99
rect 97 97 100 99
rect 39 73 40 75
rect 60 73 79 75
rect 89 73 92 75
rect 16 27 19 29
rect 39 27 51 29
rect 61 27 64 29
rect -1 -1 16 1
rect 36 -1 49 1
rect 69 -1 72 1
rect -1 -9 16 -7
rect 36 -9 49 -7
rect 69 -9 72 -7
<< polycontact >>
rect 38 344 42 348
rect -9 328 -5 332
rect 7 320 11 324
rect -10 312 -6 316
rect -9 303 -5 307
rect 38 279 42 283
rect 228 279 232 283
rect 171 253 175 257
rect 171 243 175 247
rect 335 247 339 251
rect 33 231 37 235
rect 171 233 175 237
rect 288 231 292 235
rect 304 223 308 227
rect -6 209 -2 213
rect 287 215 291 219
rect -6 197 -2 201
rect 288 206 292 210
rect 335 182 339 186
rect 35 137 39 141
rect -12 121 -8 125
rect 4 113 8 117
rect -13 105 -9 109
rect -12 96 -8 100
rect 35 72 39 76
rect 42 23 46 27
rect -5 -1 -1 3
rect -5 -9 -1 -5
<< metal1 >>
rect -9 356 70 360
rect -9 332 -5 356
rect 66 353 70 356
rect 61 349 84 353
rect -1 344 38 348
rect -10 316 -6 319
rect -1 307 3 344
rect 63 340 66 344
rect 92 340 108 344
rect 15 332 23 336
rect -5 303 3 307
rect 7 295 11 320
rect 15 320 19 332
rect 75 328 79 332
rect 63 324 79 328
rect 15 316 23 320
rect 15 303 19 316
rect 63 307 66 311
rect 75 303 79 324
rect 104 320 108 340
rect 100 316 104 320
rect 108 316 117 320
rect 15 299 23 303
rect 75 299 80 303
rect 7 291 78 295
rect 74 287 78 291
rect 63 283 82 287
rect 3 279 38 283
rect 63 274 66 278
rect 104 278 108 316
rect 228 290 232 297
rect 223 286 239 290
rect 201 278 205 282
rect 92 274 108 278
rect 59 268 63 274
rect 228 261 232 279
rect 247 278 251 282
rect 226 257 239 261
rect 260 257 268 261
rect 33 253 171 257
rect 33 242 37 253
rect 235 252 239 257
rect 226 248 231 252
rect 235 248 240 252
rect 28 238 44 242
rect 182 238 186 242
rect 6 230 10 234
rect 33 217 37 231
rect 52 230 56 234
rect 164 233 171 237
rect 227 233 231 248
rect 264 242 268 257
rect 264 233 268 238
rect 1 213 9 217
rect 33 213 41 217
rect -10 209 -6 213
rect 1 207 5 213
rect 33 207 37 213
rect 28 203 37 207
rect 164 210 168 233
rect 226 229 231 233
rect 260 229 268 233
rect 288 259 367 263
rect 288 235 292 259
rect 363 256 367 259
rect 358 252 381 256
rect 296 247 335 251
rect 287 219 291 222
rect 296 210 300 247
rect 360 243 363 247
rect 389 243 405 247
rect 312 235 320 239
rect 164 206 288 210
rect 292 206 300 210
rect -10 197 -6 201
rect 1 197 5 203
rect 1 193 9 197
rect 51 193 55 197
rect -12 149 67 153
rect -12 125 -8 149
rect 63 146 67 149
rect 58 142 81 146
rect -4 137 35 141
rect -13 109 -9 112
rect -4 100 0 137
rect 60 133 63 137
rect 89 133 105 137
rect 12 125 20 129
rect -8 96 0 100
rect 4 88 8 113
rect 12 113 16 125
rect 72 121 76 125
rect 60 117 76 121
rect 12 109 20 113
rect 12 96 16 109
rect 60 100 63 104
rect 72 96 76 117
rect 101 113 105 133
rect 97 109 101 113
rect 105 109 114 113
rect 12 92 20 96
rect 72 92 77 96
rect 4 84 75 88
rect 71 80 75 84
rect 60 76 79 80
rect 0 72 35 76
rect 60 67 63 71
rect 101 71 105 109
rect 89 67 105 71
rect 56 61 60 67
rect 164 42 168 206
rect 304 198 308 223
rect 312 223 316 235
rect 372 231 376 235
rect 360 227 376 231
rect 312 219 320 223
rect 312 206 316 219
rect 360 210 363 214
rect 372 206 376 227
rect 401 223 405 243
rect 397 219 401 223
rect 405 219 414 223
rect 312 202 320 206
rect 372 202 377 206
rect 304 194 375 198
rect 371 190 375 194
rect 360 186 379 190
rect 300 182 335 186
rect 360 177 363 181
rect 401 181 405 219
rect 389 177 405 181
rect 356 171 360 177
rect 42 38 168 42
rect 42 34 46 38
rect 37 30 53 34
rect 15 22 19 26
rect 42 6 46 23
rect 61 22 65 26
rect -7 -1 -5 3
rect 7 2 16 6
rect 42 2 49 6
rect -7 -9 -5 -5
rect 7 -10 11 2
rect 42 -2 46 2
rect 36 -6 46 -2
rect 11 -14 16 -10
rect 69 -14 73 -10
<< m2contact >>
rect -11 319 -6 324
rect 66 339 71 344
rect 75 332 80 337
rect 66 307 71 312
rect -2 279 3 284
rect 66 274 71 279
rect 166 243 171 248
rect 286 222 291 227
rect 363 242 368 247
rect 372 235 377 240
rect -14 112 -9 117
rect 63 132 68 137
rect 72 125 77 130
rect 63 100 68 105
rect -5 72 0 77
rect 63 67 68 72
rect 363 210 368 215
rect 295 182 300 187
rect 363 177 368 182
<< metal2 >>
rect 75 357 166 362
rect -6 320 3 324
rect -2 284 3 320
rect 67 312 71 339
rect 75 337 80 357
rect 67 279 71 307
rect 161 227 166 357
rect 372 260 446 265
rect 161 222 286 227
rect 291 223 300 227
rect 295 187 300 223
rect 364 215 368 242
rect 372 240 377 260
rect 364 182 368 210
rect 72 158 409 163
rect -9 113 0 117
rect -5 77 0 113
rect 64 105 68 132
rect 72 130 77 158
rect 64 72 68 100
<< labels >>
rlabel nsubstratencontact 59 264 63 268 1 vdd
rlabel metal1 95 340 96 344 7 gnd
rlabel metal1 102 316 108 320 7 gnd
rlabel polycontact -9 303 -5 307 3 A1
rlabel polycontact -10 312 -6 316 3 B1
rlabel polycontact 7 320 11 324 1 B1_bar
rlabel polycontact -9 328 -5 332 3 A1_bar
rlabel metal1 178 238 179 241 3 vdd
rlabel metal1 169 233 170 236 3 G0
rlabel m2contact 169 243 170 246 3 P1
rlabel metal1 169 253 170 256 3 G1
rlabel metal1 202 278 203 282 7 vdd
rlabel metal1 250 278 251 282 7 gnd
rlabel metal1 230 265 231 270 7 C2_bar
rlabel metal1 229 296 231 297 5 C2
rlabel metal1 265 229 266 232 8 gnd
rlabel nsubstratencontact 356 167 360 171 1 vdd
rlabel metal1 392 243 393 247 7 gnd
rlabel metal1 399 219 405 223 7 gnd
rlabel metal1 99 109 105 113 7 gnd
rlabel nsubstratencontact 56 57 60 61 1 vdd
rlabel polycontact -12 96 -8 100 3 A0
rlabel polycontact -13 105 -9 109 3 B0
rlabel polycontact -12 121 -8 125 3 A0_bar
rlabel metal1 92 133 93 137 7 gnd
rlabel metal2 73 161 76 162 1 S0
rlabel metal2 373 261 376 263 1 S1
rlabel polycontact 287 215 291 219 1 P1
rlabel polycontact 288 206 292 210 1 G0
rlabel polycontact 304 223 308 227 1 P1_bar
rlabel polycontact 288 231 292 235 1 G0_bar
rlabel metal1 34 248 36 249 1 G1
rlabel metal1 35 220 36 225 1 G1_bar
rlabel metal1 -10 210 -9 212 3 B1
rlabel metal1 -10 198 -9 200 3 A1
rlabel metal1 53 193 55 194 8 gnd
rlabel metal1 1 193 2 197 3 vdd
rlabel metal1 7 230 8 234 7 vdd
rlabel metal1 55 230 56 234 7 gnd
rlabel psubstratepcontact 73 -14 77 -10 7 gnd
rlabel nsubstratencontact 7 -14 11 -10 7 vdd
rlabel metal1 -7 -9 -5 -7 3 A0
rlabel metal1 -7 -1 -5 1 3 B0
rlabel metal1 42 13 46 15 1 G0_bar
rlabel metal1 64 22 65 26 7 gnd
rlabel metal1 16 22 17 26 7 vdd
rlabel metal1 43 40 45 41 1 G0
<< end >>
