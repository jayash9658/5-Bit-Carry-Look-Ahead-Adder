magic
tech scmos
timestamp 1764679931
<< nwell >>
rect -119 896 -87 984
rect 37 980 85 1001
rect 28 923 85 980
rect 286 952 323 983
rect 43 904 85 923
rect 63 899 85 904
rect -119 799 -87 887
rect 10 860 47 887
rect 9 857 47 860
rect 9 821 46 857
rect 262 836 320 952
rect 424 912 456 1000
rect 432 847 480 868
rect 579 857 611 945
rect -119 700 -87 788
rect 37 785 85 806
rect 423 790 480 847
rect 28 728 85 785
rect 286 742 323 773
rect 438 766 480 790
rect 43 709 85 728
rect 63 704 85 709
rect -119 601 -87 689
rect 10 660 47 687
rect 9 657 47 660
rect 9 621 46 657
rect 262 646 320 742
rect 432 653 480 674
rect 579 663 611 751
rect -119 503 -87 591
rect 37 587 85 608
rect 423 596 480 653
rect 28 530 85 587
rect 438 572 480 596
rect 43 511 85 530
rect 63 506 85 511
rect 261 521 324 552
rect -119 405 -87 493
rect 10 466 47 493
rect 9 463 47 466
rect 9 427 46 463
rect 261 454 323 521
rect 432 440 480 461
rect 579 450 611 538
rect -119 306 -87 394
rect 37 389 85 410
rect 28 332 85 389
rect 423 383 480 440
rect 438 359 480 383
rect 43 308 85 332
rect 287 316 324 347
rect 260 313 324 316
rect -119 208 -87 296
rect 10 269 47 296
rect 260 269 325 313
rect 432 286 480 307
rect 579 296 611 384
rect 9 266 47 269
rect 9 230 46 266
rect 423 229 480 286
rect -119 111 -87 199
rect 37 186 85 207
rect 438 205 480 229
rect 579 188 611 276
rect 28 129 85 186
rect 43 110 85 129
rect 63 105 85 110
rect -119 11 -87 99
rect 10 54 47 81
rect 9 51 47 54
rect 9 15 46 51
<< ntransistor >>
rect 468 987 478 989
rect 93 983 103 985
rect -75 971 -65 973
rect 91 967 111 969
rect 468 971 478 973
rect 329 965 339 967
rect 91 959 111 961
rect 468 963 478 965
rect -75 955 -65 957
rect 91 951 111 953
rect -75 947 -65 949
rect 468 947 478 949
rect 91 942 111 944
rect 328 939 348 941
rect -75 931 -65 933
rect 468 939 478 941
rect 328 929 348 931
rect 623 932 633 934
rect -75 923 -65 925
rect 468 923 478 925
rect 93 918 103 920
rect 623 916 633 918
rect 328 913 348 915
rect -75 907 -65 909
rect 623 908 633 910
rect 328 903 348 905
rect 328 893 348 895
rect 623 892 633 894
rect 328 883 348 885
rect 623 884 633 886
rect -75 874 -65 876
rect 53 869 63 871
rect 328 867 348 869
rect 623 868 633 870
rect -75 858 -65 860
rect 328 857 348 859
rect -75 850 -65 852
rect 488 850 498 852
rect 328 847 348 849
rect 52 844 62 846
rect -75 834 -65 836
rect 52 832 62 834
rect 486 834 506 836
rect -75 826 -65 828
rect 486 826 506 828
rect 486 818 506 820
rect -75 810 -65 812
rect 486 809 506 811
rect 93 788 103 790
rect 488 785 498 787
rect -75 775 -65 777
rect 91 772 111 774
rect 91 764 111 766
rect -75 759 -65 761
rect 91 756 111 758
rect -75 751 -65 753
rect 329 755 339 757
rect 91 747 111 749
rect 623 738 633 740
rect -75 735 -65 737
rect -75 727 -65 729
rect 328 729 348 731
rect 93 723 103 725
rect 623 722 633 724
rect 328 719 348 721
rect -75 711 -65 713
rect 623 714 633 716
rect 328 709 348 711
rect 623 698 633 700
rect 328 693 348 695
rect 623 690 633 692
rect 328 683 348 685
rect -75 676 -65 678
rect 53 669 63 671
rect 623 674 633 676
rect 328 667 348 669
rect -75 660 -65 662
rect 328 657 348 659
rect -75 652 -65 654
rect 488 656 498 658
rect 52 644 62 646
rect -75 636 -65 638
rect 486 640 506 642
rect 52 632 62 634
rect -75 628 -65 630
rect 486 632 506 634
rect 486 624 506 626
rect 486 615 506 617
rect -75 612 -65 614
rect 93 590 103 592
rect 488 591 498 593
rect -75 578 -65 580
rect 91 574 111 576
rect 91 566 111 568
rect -75 562 -65 564
rect 91 558 111 560
rect -75 554 -65 556
rect 91 549 111 551
rect -75 538 -65 540
rect 330 534 340 536
rect -75 530 -65 532
rect 93 525 103 527
rect 623 525 633 527
rect -75 514 -65 516
rect 330 509 350 511
rect 623 509 633 511
rect 330 501 350 503
rect 623 501 633 503
rect 330 485 350 487
rect -75 480 -65 482
rect 53 475 63 477
rect 623 485 633 487
rect 330 475 350 477
rect 623 477 633 479
rect -75 464 -65 466
rect 330 465 350 467
rect 623 461 633 463
rect -75 456 -65 458
rect 52 450 62 452
rect -75 440 -65 442
rect 488 443 498 445
rect 52 438 62 440
rect -75 432 -65 434
rect 486 427 506 429
rect 486 419 506 421
rect -75 416 -65 418
rect 486 411 506 413
rect 486 402 506 404
rect 93 392 103 394
rect -75 381 -65 383
rect 91 376 111 378
rect 488 378 498 380
rect -75 365 -65 367
rect 623 371 633 373
rect 91 368 111 370
rect 91 360 111 362
rect -75 357 -65 359
rect 623 355 633 357
rect 91 351 111 353
rect 623 347 633 349
rect -75 341 -65 343
rect -75 333 -65 335
rect 330 329 340 331
rect 623 331 633 333
rect 93 327 103 329
rect 623 323 633 325
rect -75 317 -65 319
rect 623 307 633 309
rect 333 300 353 302
rect 333 290 353 292
rect -75 283 -65 285
rect 53 278 63 280
rect 488 289 498 291
rect 333 280 353 282
rect 486 273 506 275
rect -75 267 -65 269
rect 486 265 506 267
rect -75 259 -65 261
rect 623 263 633 265
rect 486 257 506 259
rect 52 253 62 255
rect -75 243 -65 245
rect 486 248 506 250
rect 623 247 633 249
rect 52 241 62 243
rect -75 235 -65 237
rect 623 239 633 241
rect 488 224 498 226
rect -75 219 -65 221
rect 623 223 633 225
rect 623 215 633 217
rect 623 199 633 201
rect 93 189 103 191
rect -75 186 -65 188
rect -75 170 -65 172
rect 91 173 111 175
rect 91 165 111 167
rect -75 162 -65 164
rect 91 157 111 159
rect -75 146 -65 148
rect 91 148 111 150
rect -75 138 -65 140
rect -75 122 -65 124
rect 93 124 103 126
rect -75 86 -65 88
rect -75 70 -65 72
rect -75 62 -65 64
rect 53 63 63 65
rect -75 46 -65 48
rect -75 38 -65 40
rect 52 38 62 40
rect 52 26 62 28
rect -75 22 -65 24
<< ptransistor >>
rect 430 987 450 989
rect 54 983 74 985
rect -113 971 -93 973
rect 34 967 74 969
rect 297 965 317 967
rect 34 959 74 961
rect 430 963 450 965
rect 34 951 74 953
rect -113 947 -93 949
rect 430 947 450 949
rect 34 942 74 944
rect 274 939 314 941
rect -113 931 -93 933
rect 274 929 314 931
rect 430 931 450 933
rect 585 932 605 934
rect 430 923 450 925
rect 54 918 74 920
rect -113 915 -93 917
rect 274 913 314 915
rect -113 907 -93 909
rect 585 908 605 910
rect 274 903 314 905
rect 274 893 314 895
rect 585 892 605 894
rect 274 883 314 885
rect -113 874 -93 876
rect 585 876 605 878
rect 21 869 41 871
rect 274 867 314 869
rect 585 868 605 870
rect 274 857 314 859
rect -113 850 -93 852
rect 449 850 469 852
rect 274 847 314 849
rect 20 844 40 846
rect -113 834 -93 836
rect 20 832 40 834
rect 429 834 469 836
rect 429 826 469 828
rect -113 818 -93 820
rect 429 818 469 820
rect -113 810 -93 812
rect 429 809 469 811
rect 54 788 74 790
rect 449 785 469 787
rect -113 775 -93 777
rect 34 772 74 774
rect 34 764 74 766
rect 34 756 74 758
rect -113 751 -93 753
rect 297 755 317 757
rect 34 747 74 749
rect 585 738 605 740
rect -113 735 -93 737
rect 274 729 314 731
rect 54 723 74 725
rect -113 719 -93 721
rect 274 719 314 721
rect -113 711 -93 713
rect 585 714 605 716
rect 274 709 314 711
rect 585 698 605 700
rect 274 693 314 695
rect 274 683 314 685
rect 585 682 605 684
rect -113 676 -93 678
rect 21 669 41 671
rect 585 674 605 676
rect 274 667 314 669
rect 274 657 314 659
rect -113 652 -93 654
rect 449 656 469 658
rect 20 644 40 646
rect -113 636 -93 638
rect 429 640 469 642
rect 20 632 40 634
rect 429 632 469 634
rect 429 624 469 626
rect -113 620 -93 622
rect 429 615 469 617
rect -113 612 -93 614
rect 54 590 74 592
rect 449 591 469 593
rect -113 578 -93 580
rect 34 574 74 576
rect 34 566 74 568
rect 34 558 74 560
rect -113 554 -93 556
rect 34 549 74 551
rect -113 538 -93 540
rect 298 534 318 536
rect 54 525 74 527
rect 585 525 605 527
rect -113 522 -93 524
rect -113 514 -93 516
rect 276 509 316 511
rect 276 501 316 503
rect 585 501 605 503
rect 276 485 316 487
rect -113 480 -93 482
rect 21 475 41 477
rect 585 485 605 487
rect 276 475 316 477
rect 585 469 605 471
rect 276 465 316 467
rect 585 461 605 463
rect -113 456 -93 458
rect 20 450 40 452
rect -113 440 -93 442
rect 449 443 469 445
rect 20 438 40 440
rect 429 427 469 429
rect -113 424 -93 426
rect 429 419 469 421
rect -113 416 -93 418
rect 429 411 469 413
rect 429 402 469 404
rect 54 392 74 394
rect -113 381 -93 383
rect 34 376 74 378
rect 449 378 469 380
rect 585 371 605 373
rect 34 368 74 370
rect 34 360 74 362
rect -113 357 -93 359
rect 34 351 74 353
rect 585 347 605 349
rect -113 341 -93 343
rect -113 325 -93 327
rect 298 329 318 331
rect 585 331 605 333
rect 54 327 74 329
rect -113 317 -93 319
rect 585 315 605 317
rect 585 307 605 309
rect 279 300 319 302
rect 279 290 319 292
rect -113 283 -93 285
rect 21 278 41 280
rect 449 289 469 291
rect 279 280 319 282
rect 429 273 469 275
rect 429 265 469 267
rect -113 259 -93 261
rect 585 263 605 265
rect 429 257 469 259
rect 20 253 40 255
rect -113 243 -93 245
rect 429 248 469 250
rect 20 241 40 243
rect 585 239 605 241
rect -113 227 -93 229
rect 449 224 469 226
rect -113 219 -93 221
rect 585 223 605 225
rect 585 207 605 209
rect 585 199 605 201
rect 54 189 74 191
rect -113 186 -93 188
rect 34 173 74 175
rect 34 165 74 167
rect -113 162 -93 164
rect 34 157 74 159
rect -113 146 -93 148
rect 34 148 74 150
rect -113 130 -93 132
rect -113 122 -93 124
rect 54 124 74 126
rect -113 86 -93 88
rect -113 62 -93 64
rect 21 63 41 65
rect -113 46 -93 48
rect 20 38 40 40
rect -113 30 -93 32
rect 20 26 40 28
rect -113 22 -93 24
<< ndiffusion >>
rect 93 987 95 991
rect 99 987 103 991
rect 472 990 478 994
rect 468 989 478 990
rect 93 985 103 987
rect 93 982 103 983
rect 468 986 478 987
rect 468 982 474 986
rect 93 978 99 982
rect -71 974 -65 978
rect 472 974 478 978
rect -75 973 -65 974
rect -75 970 -65 971
rect -75 966 -69 970
rect 95 970 111 974
rect 468 973 478 974
rect 91 969 111 970
rect 329 968 331 972
rect 335 968 339 972
rect 329 967 339 968
rect -71 958 -65 962
rect 91 961 111 967
rect 468 965 478 971
rect 329 964 339 965
rect 329 960 335 964
rect -75 957 -65 958
rect -75 949 -65 955
rect 91 958 111 959
rect 468 962 478 963
rect 468 958 474 962
rect 91 954 107 958
rect 91 953 111 954
rect -75 946 -65 947
rect -75 942 -69 946
rect 91 944 111 951
rect 468 950 474 954
rect 468 949 478 950
rect -75 934 -69 938
rect 91 941 111 942
rect 95 937 111 941
rect 332 942 348 946
rect 328 941 348 942
rect -75 933 -65 934
rect -75 925 -65 931
rect 328 937 348 939
rect 468 941 478 947
rect 468 938 478 939
rect 328 933 344 937
rect 472 934 478 938
rect 627 935 633 939
rect 623 934 633 935
rect 328 931 348 933
rect -75 922 -65 923
rect -71 918 -65 922
rect 97 921 103 925
rect 328 928 348 929
rect 328 924 344 928
rect 472 926 478 930
rect 623 931 633 932
rect 623 927 629 931
rect 468 925 478 926
rect 93 920 103 921
rect -71 910 -65 914
rect 93 916 103 918
rect 93 912 99 916
rect 332 916 348 920
rect 468 922 478 923
rect 468 918 474 922
rect 627 919 633 923
rect 623 918 633 919
rect 328 915 348 916
rect -75 909 -65 910
rect -75 906 -65 907
rect -75 902 -69 906
rect 328 911 348 913
rect 328 907 344 911
rect 623 910 633 916
rect 328 905 348 907
rect 623 907 633 908
rect 623 903 629 907
rect 328 901 348 903
rect 332 897 348 901
rect 328 895 348 897
rect 328 891 348 893
rect 623 895 629 899
rect 623 894 633 895
rect 328 887 344 891
rect 328 885 348 887
rect 623 886 633 892
rect 623 883 633 884
rect -71 877 -65 881
rect 328 882 348 883
rect 328 878 344 882
rect 627 879 633 883
rect -75 876 -65 877
rect -75 873 -65 874
rect -75 869 -69 873
rect 53 872 55 876
rect 59 872 63 876
rect 53 871 63 872
rect -71 861 -65 865
rect 53 868 63 869
rect 53 864 59 868
rect 332 870 348 874
rect 328 869 348 870
rect 627 871 633 875
rect 623 870 633 871
rect -75 860 -65 861
rect -75 852 -65 858
rect 328 865 348 867
rect 328 861 344 865
rect 623 867 633 868
rect 623 863 629 867
rect 328 859 348 861
rect -75 849 -65 850
rect -75 845 -69 849
rect 56 847 62 851
rect 52 846 62 847
rect 328 849 348 857
rect 488 854 490 858
rect 494 854 498 858
rect 488 852 498 854
rect -75 837 -69 841
rect -75 836 -65 837
rect -75 828 -65 834
rect 52 834 62 844
rect 328 846 348 847
rect 328 842 344 846
rect 488 849 498 850
rect 488 845 494 849
rect 490 837 506 841
rect 486 836 506 837
rect 52 831 62 832
rect 52 827 58 831
rect -75 825 -65 826
rect 486 828 506 834
rect -71 821 -65 825
rect 486 825 506 826
rect 486 821 502 825
rect 486 820 506 821
rect -71 813 -65 817
rect -75 812 -65 813
rect -75 809 -65 810
rect -75 805 -69 809
rect 486 811 506 818
rect 486 808 506 809
rect 490 804 506 808
rect 93 792 95 796
rect 99 792 103 796
rect 93 790 103 792
rect 93 787 103 788
rect 93 783 99 787
rect 492 788 498 792
rect 488 787 498 788
rect -71 778 -65 782
rect 488 783 498 785
rect 488 779 494 783
rect -75 777 -65 778
rect -75 774 -65 775
rect -75 770 -69 774
rect 95 775 111 779
rect 91 774 111 775
rect -71 762 -65 766
rect 91 766 111 772
rect -75 761 -65 762
rect -75 753 -65 759
rect 91 763 111 764
rect 91 759 107 763
rect 91 758 111 759
rect 329 758 331 762
rect 335 758 339 762
rect 329 757 339 758
rect -75 750 -65 751
rect -75 746 -69 750
rect 91 749 111 756
rect 329 754 339 755
rect 329 750 335 754
rect 91 746 111 747
rect 95 742 111 746
rect -75 738 -69 742
rect 627 741 633 745
rect 623 740 633 741
rect -75 737 -65 738
rect -75 729 -65 735
rect -75 726 -65 727
rect -71 722 -65 726
rect 97 726 103 730
rect 332 732 348 736
rect 623 737 633 738
rect 623 733 629 737
rect 328 731 348 732
rect 93 725 103 726
rect -71 714 -65 718
rect 93 721 103 723
rect 93 717 99 721
rect 328 727 348 729
rect 328 723 344 727
rect 627 725 633 729
rect 623 724 633 725
rect 328 721 348 723
rect -75 713 -65 714
rect -75 710 -65 711
rect -75 706 -69 710
rect 328 711 348 719
rect 623 716 633 722
rect 623 713 633 714
rect 623 709 629 713
rect 328 708 348 709
rect 332 704 348 708
rect 332 696 348 700
rect 623 701 629 705
rect 623 700 633 701
rect 328 695 348 696
rect -71 679 -65 683
rect 328 691 348 693
rect 332 687 348 691
rect 623 692 633 698
rect 623 689 633 690
rect 328 685 348 687
rect 627 685 633 689
rect -75 678 -65 679
rect 328 682 348 683
rect 328 678 344 682
rect -75 675 -65 676
rect -75 671 -69 675
rect 53 672 55 676
rect 59 672 63 676
rect 53 671 63 672
rect -71 663 -65 667
rect 53 668 63 669
rect 53 664 59 668
rect 332 670 348 674
rect 627 677 633 681
rect 623 676 633 677
rect 328 669 348 670
rect 623 673 633 674
rect 623 669 629 673
rect -75 662 -65 663
rect -75 654 -65 660
rect 328 665 348 667
rect 332 661 348 665
rect 328 659 348 661
rect 328 656 348 657
rect 328 652 344 656
rect 488 660 490 664
rect 494 660 498 664
rect 488 658 498 660
rect -75 651 -65 652
rect 488 655 498 656
rect 488 651 494 655
rect -75 647 -69 651
rect 56 647 62 651
rect 52 646 62 647
rect -75 639 -69 643
rect -75 638 -65 639
rect -75 630 -65 636
rect 52 634 62 644
rect 490 643 506 647
rect 486 642 506 643
rect -75 627 -65 628
rect 52 631 62 632
rect 486 634 506 640
rect 52 627 58 631
rect -71 623 -65 627
rect 486 631 506 632
rect 486 627 502 631
rect 486 626 506 627
rect -71 615 -65 619
rect -75 614 -65 615
rect 486 617 506 624
rect -75 611 -65 612
rect -75 607 -69 611
rect 486 614 506 615
rect 490 610 506 614
rect 93 594 95 598
rect 99 594 103 598
rect 93 592 103 594
rect 492 594 498 598
rect 488 593 498 594
rect 93 589 103 590
rect 93 585 99 589
rect 488 589 498 591
rect 488 585 494 589
rect -71 581 -65 585
rect -75 580 -65 581
rect -75 577 -65 578
rect -75 573 -69 577
rect 95 577 111 581
rect 91 576 111 577
rect -71 565 -65 569
rect 91 568 111 574
rect -75 564 -65 565
rect -75 556 -65 562
rect 91 565 111 566
rect 91 561 107 565
rect 91 560 111 561
rect -75 553 -65 554
rect -75 549 -69 553
rect 91 551 111 558
rect -75 541 -69 545
rect 91 548 111 549
rect 95 544 111 548
rect -75 540 -65 541
rect -75 532 -65 538
rect 330 537 332 541
rect 336 537 340 541
rect 330 536 340 537
rect -75 529 -65 530
rect -71 525 -65 529
rect 97 528 103 532
rect 330 533 340 534
rect 330 529 336 533
rect 93 527 103 528
rect 627 528 633 532
rect 623 527 633 528
rect -71 517 -65 521
rect 93 523 103 525
rect 93 519 99 523
rect 623 524 633 525
rect 623 520 629 524
rect -75 516 -65 517
rect -75 513 -65 514
rect -75 509 -69 513
rect 334 512 350 516
rect 627 512 633 516
rect 330 511 350 512
rect 623 511 633 512
rect 330 508 350 509
rect 330 504 346 508
rect 330 503 350 504
rect 623 503 633 509
rect 330 500 350 501
rect 330 496 346 500
rect 623 500 633 501
rect 623 496 629 500
rect -71 483 -65 487
rect 330 488 346 492
rect 330 487 350 488
rect -75 482 -65 483
rect -75 479 -65 480
rect -75 475 -69 479
rect 53 478 55 482
rect 59 478 63 482
rect 53 477 63 478
rect -71 467 -65 471
rect 53 474 63 475
rect 330 483 350 485
rect 623 488 629 492
rect 623 487 633 488
rect 334 479 350 483
rect 330 477 350 479
rect 623 479 633 485
rect 623 476 633 477
rect 53 470 59 474
rect -75 466 -65 467
rect -75 458 -65 464
rect 330 473 350 475
rect 334 469 350 473
rect 627 472 633 476
rect 330 467 350 469
rect 330 464 350 465
rect 330 460 346 464
rect 627 464 633 468
rect 623 463 633 464
rect -75 455 -65 456
rect -75 451 -69 455
rect 56 453 62 457
rect 623 460 633 461
rect 623 456 629 460
rect 52 452 62 453
rect -75 443 -69 447
rect -75 442 -65 443
rect -75 434 -65 440
rect 52 440 62 450
rect 488 447 490 451
rect 494 447 498 451
rect 488 445 498 447
rect 488 442 498 443
rect 488 438 494 442
rect 52 437 62 438
rect 52 433 58 437
rect -75 431 -65 432
rect -71 427 -65 431
rect 490 430 506 434
rect 486 429 506 430
rect -71 419 -65 423
rect -75 418 -65 419
rect 486 421 506 427
rect -75 415 -65 416
rect -75 411 -69 415
rect 486 418 506 419
rect 486 414 502 418
rect 486 413 506 414
rect 486 404 506 411
rect 93 396 95 400
rect 99 396 103 400
rect 486 401 506 402
rect 490 397 506 401
rect 93 394 103 396
rect -71 384 -65 388
rect 93 391 103 392
rect 93 387 99 391
rect -75 383 -65 384
rect -75 380 -65 381
rect -75 376 -69 380
rect 95 379 111 383
rect 91 378 111 379
rect 492 381 498 385
rect 488 380 498 381
rect -71 368 -65 372
rect -75 367 -65 368
rect -75 359 -65 365
rect 91 370 111 376
rect 488 376 498 378
rect 488 372 494 376
rect 627 374 633 378
rect 623 373 633 374
rect 91 367 111 368
rect 91 363 107 367
rect 623 370 633 371
rect 623 366 629 370
rect 91 362 111 363
rect -75 356 -65 357
rect -75 352 -69 356
rect 91 353 111 360
rect 627 358 633 362
rect 623 357 633 358
rect -75 344 -69 348
rect 91 350 111 351
rect 95 346 111 350
rect 623 349 633 355
rect -75 343 -65 344
rect -75 335 -65 341
rect 623 346 633 347
rect 623 342 629 346
rect -75 332 -65 333
rect -71 328 -65 332
rect 97 330 103 334
rect 330 332 332 336
rect 336 332 340 336
rect 330 331 340 332
rect 93 329 103 330
rect 623 334 629 338
rect 623 333 633 334
rect -71 320 -65 324
rect 93 325 103 327
rect 93 321 99 325
rect 330 328 340 329
rect 330 324 336 328
rect 623 325 633 331
rect 623 322 633 323
rect -75 319 -65 320
rect 627 318 633 322
rect -75 316 -65 317
rect -75 312 -69 316
rect 333 303 349 307
rect 627 310 633 314
rect 623 309 633 310
rect 333 302 353 303
rect 623 306 633 307
rect 623 302 629 306
rect -71 286 -65 290
rect 333 298 353 300
rect 337 294 353 298
rect 333 292 353 294
rect -75 285 -65 286
rect -75 282 -65 283
rect -75 278 -69 282
rect 53 281 55 285
rect 59 281 63 285
rect 53 280 63 281
rect 333 282 353 290
rect 488 293 490 297
rect 494 293 498 297
rect 488 291 498 293
rect 488 288 498 289
rect 488 284 494 288
rect -71 270 -65 274
rect 53 277 63 278
rect 53 273 59 277
rect 333 279 353 280
rect 333 275 349 279
rect 490 276 506 280
rect 486 275 506 276
rect -75 269 -65 270
rect -75 261 -65 267
rect 486 267 506 273
rect 627 266 633 270
rect 623 265 633 266
rect -75 258 -65 259
rect -75 254 -69 258
rect 56 256 62 260
rect 486 264 506 265
rect 486 260 502 264
rect 486 259 506 260
rect 623 262 633 263
rect 623 258 629 262
rect 52 255 62 256
rect -75 246 -69 250
rect -75 245 -65 246
rect -75 237 -65 243
rect 52 243 62 253
rect 486 250 506 257
rect 627 250 633 254
rect 623 249 633 250
rect 486 247 506 248
rect 490 243 506 247
rect 623 241 633 247
rect 52 240 62 241
rect 52 236 58 240
rect -75 234 -65 235
rect 623 238 633 239
rect 623 234 629 238
rect -71 230 -65 234
rect -71 222 -65 226
rect 492 227 498 231
rect 488 226 498 227
rect -75 221 -65 222
rect -75 218 -65 219
rect 488 222 498 224
rect 623 226 629 230
rect 623 225 633 226
rect 488 218 494 222
rect -75 214 -69 218
rect 623 217 633 223
rect 623 214 633 215
rect 627 210 633 214
rect 627 202 633 206
rect 623 201 633 202
rect -71 189 -65 193
rect -75 188 -65 189
rect 93 193 95 197
rect 99 193 103 197
rect 623 198 633 199
rect 623 194 629 198
rect 93 191 103 193
rect -75 185 -65 186
rect -75 181 -69 185
rect 93 188 103 189
rect 93 184 99 188
rect -71 173 -65 177
rect -75 172 -65 173
rect -75 164 -65 170
rect 95 176 111 180
rect 91 175 111 176
rect 91 167 111 173
rect -75 161 -65 162
rect -75 157 -69 161
rect 91 164 111 165
rect 91 160 107 164
rect 91 159 111 160
rect -75 149 -69 153
rect -75 148 -65 149
rect -75 140 -65 146
rect 91 150 111 157
rect 91 147 111 148
rect 95 143 111 147
rect -75 137 -65 138
rect -71 133 -65 137
rect -71 125 -65 129
rect -75 124 -65 125
rect 97 127 103 131
rect 93 126 103 127
rect -75 121 -65 122
rect -75 117 -69 121
rect 93 122 103 124
rect 93 118 99 122
rect -71 89 -65 93
rect -75 88 -65 89
rect -75 85 -65 86
rect -75 81 -69 85
rect -71 73 -65 77
rect -75 72 -65 73
rect -75 64 -65 70
rect 53 66 55 70
rect 59 66 63 70
rect 53 65 63 66
rect -75 61 -65 62
rect -75 57 -69 61
rect 53 62 63 63
rect 53 58 59 62
rect -75 49 -69 53
rect -75 48 -65 49
rect -75 40 -65 46
rect -75 37 -65 38
rect 56 41 62 45
rect 52 40 62 41
rect -71 33 -65 37
rect -71 25 -65 29
rect 52 28 62 38
rect -75 24 -65 25
rect -75 21 -65 22
rect 52 25 62 26
rect 52 21 58 25
rect -75 17 -69 21
<< pdiffusion >>
rect 54 987 68 991
rect 72 987 74 991
rect 54 985 74 987
rect 430 990 446 994
rect 430 989 450 990
rect 430 986 450 987
rect 54 982 74 983
rect 54 978 70 982
rect 434 982 450 986
rect -113 974 -97 978
rect -113 973 -93 974
rect 54 977 74 978
rect -113 970 -93 971
rect -109 966 -93 970
rect 38 970 74 974
rect 34 969 74 970
rect 297 968 311 972
rect 315 968 317 972
rect 297 967 317 968
rect 34 966 74 967
rect 34 962 70 966
rect 34 961 74 962
rect 430 966 446 970
rect 430 965 450 966
rect 297 964 317 965
rect 301 960 317 964
rect 430 962 450 963
rect 34 958 74 959
rect -113 950 -97 954
rect -113 949 -93 950
rect 38 954 74 958
rect 34 953 74 954
rect 434 958 450 962
rect 34 949 74 951
rect -113 946 -93 947
rect -109 942 -93 946
rect 34 945 70 949
rect 34 944 74 945
rect 430 950 446 954
rect 430 949 450 950
rect 430 946 450 947
rect 274 942 310 946
rect 34 941 74 942
rect -113 934 -97 938
rect -113 933 -93 934
rect 38 937 74 941
rect 274 941 314 942
rect 434 942 450 946
rect 274 937 314 939
rect -113 930 -93 931
rect -109 926 -93 930
rect 278 933 314 937
rect 274 931 314 933
rect 430 934 446 938
rect 585 935 601 939
rect 585 934 605 935
rect 430 933 450 934
rect 585 931 605 932
rect 274 928 314 929
rect 54 925 74 926
rect -113 918 -97 922
rect 54 921 70 925
rect -113 917 -93 918
rect 54 920 74 921
rect 274 924 310 928
rect 430 925 450 931
rect 589 927 605 931
rect 430 922 450 923
rect 54 916 74 918
rect -113 909 -93 915
rect 54 912 70 916
rect 278 916 314 920
rect 274 915 314 916
rect 434 918 450 922
rect 274 911 314 913
rect 278 907 314 911
rect -113 906 -93 907
rect -109 902 -93 906
rect 274 905 314 907
rect 585 911 601 915
rect 585 910 605 911
rect 585 907 605 908
rect 589 903 605 907
rect 274 901 314 903
rect 274 897 310 901
rect 274 895 314 897
rect 585 895 601 899
rect 274 891 314 893
rect 278 887 314 891
rect 274 885 314 887
rect 585 894 605 895
rect 585 891 605 892
rect 589 887 605 891
rect 274 882 314 883
rect -113 877 -97 881
rect -113 876 -93 877
rect 274 878 310 882
rect 585 879 601 883
rect -113 873 -93 874
rect -109 869 -93 873
rect 21 872 35 876
rect 39 872 41 876
rect 21 871 41 872
rect 585 878 605 879
rect 278 870 314 874
rect 21 868 41 869
rect 25 864 41 868
rect 274 869 314 870
rect 585 870 605 876
rect 585 867 605 868
rect 274 865 314 867
rect 278 861 314 865
rect -113 853 -97 857
rect -113 852 -93 853
rect 274 859 314 861
rect 589 863 605 867
rect 274 855 314 857
rect 274 851 310 855
rect -113 849 -93 850
rect -109 845 -93 849
rect 24 847 40 851
rect 20 846 40 847
rect 274 849 314 851
rect 449 854 463 858
rect 467 854 469 858
rect 449 852 469 854
rect 449 849 469 850
rect 274 846 314 847
rect 20 841 40 844
rect -113 837 -97 841
rect -113 836 -93 837
rect 20 837 35 841
rect 39 837 40 841
rect -113 833 -93 834
rect -109 829 -93 833
rect 20 834 40 837
rect 278 842 314 846
rect 449 845 465 849
rect 449 844 469 845
rect 433 837 469 841
rect 429 836 469 837
rect 429 833 469 834
rect 20 831 40 832
rect 24 827 40 831
rect 429 829 465 833
rect 429 828 469 829
rect 429 825 469 826
rect -113 821 -97 825
rect 433 821 469 825
rect -113 820 -93 821
rect -113 812 -93 818
rect 429 820 469 821
rect 429 816 469 818
rect 429 812 465 816
rect -113 809 -93 810
rect -109 805 -93 809
rect 429 811 469 812
rect 429 808 469 809
rect 433 804 469 808
rect 54 792 68 796
rect 72 792 74 796
rect 54 790 74 792
rect 449 792 469 793
rect 449 788 465 792
rect 54 787 74 788
rect 54 783 70 787
rect 449 787 469 788
rect 449 783 469 785
rect 54 782 74 783
rect -113 778 -97 782
rect -113 777 -93 778
rect 449 779 465 783
rect 38 775 74 779
rect -113 774 -93 775
rect -109 770 -93 774
rect 34 774 74 775
rect 34 771 74 772
rect 34 767 70 771
rect 34 766 74 767
rect 34 763 74 764
rect -113 754 -97 758
rect -113 753 -93 754
rect 38 759 74 763
rect 34 758 74 759
rect 297 758 311 762
rect 315 758 317 762
rect 297 757 317 758
rect 34 754 74 756
rect -113 750 -93 751
rect -109 746 -93 750
rect 34 750 70 754
rect 34 749 74 750
rect 297 754 317 755
rect 301 750 317 754
rect 34 746 74 747
rect 38 742 74 746
rect -113 738 -97 742
rect -113 737 -93 738
rect 585 741 601 745
rect 585 740 605 741
rect -113 734 -93 735
rect -109 730 -93 734
rect 585 737 605 738
rect 278 732 314 736
rect 54 730 74 731
rect 54 726 70 730
rect -113 722 -97 726
rect 54 725 74 726
rect 274 731 314 732
rect 589 733 605 737
rect 274 727 314 729
rect 278 723 314 727
rect -113 721 -93 722
rect 54 721 74 723
rect -113 713 -93 719
rect 54 717 70 721
rect 274 721 314 723
rect 274 717 314 719
rect 274 713 310 717
rect -113 710 -93 711
rect -109 706 -93 710
rect 274 711 314 713
rect 585 717 601 721
rect 585 716 605 717
rect 585 713 605 714
rect 589 709 605 713
rect 274 708 314 709
rect 278 704 314 708
rect 585 701 601 705
rect 274 696 310 700
rect 274 695 314 696
rect 585 700 605 701
rect 585 697 605 698
rect 589 693 605 697
rect 274 691 314 693
rect 278 687 314 691
rect -113 679 -97 683
rect -113 678 -93 679
rect 274 685 314 687
rect 585 685 601 689
rect 274 682 314 683
rect 278 678 314 682
rect 585 684 605 685
rect -113 675 -93 676
rect -109 671 -93 675
rect 21 672 35 676
rect 39 672 41 676
rect 21 671 41 672
rect 274 670 310 674
rect 21 668 41 669
rect 25 664 41 668
rect 274 669 314 670
rect 585 676 605 682
rect 585 673 605 674
rect 589 669 605 673
rect 274 665 314 667
rect -113 655 -97 659
rect -113 654 -93 655
rect 278 661 314 665
rect 274 659 314 661
rect 449 660 463 664
rect 467 660 469 664
rect 274 656 314 657
rect 278 652 314 656
rect 449 658 469 660
rect 449 655 469 656
rect -113 651 -93 652
rect -109 647 -93 651
rect 449 651 465 655
rect 24 647 40 651
rect 20 646 40 647
rect 449 650 469 651
rect -113 639 -97 643
rect -113 638 -93 639
rect 20 641 40 644
rect -113 635 -93 636
rect -109 631 -93 635
rect 20 637 35 641
rect 39 637 40 641
rect 20 634 40 637
rect 433 643 469 647
rect 429 642 469 643
rect 429 639 469 640
rect 429 635 465 639
rect 20 631 40 632
rect 24 627 40 631
rect 429 634 469 635
rect 429 631 469 632
rect 433 627 469 631
rect -113 623 -97 627
rect 429 626 469 627
rect -113 622 -93 623
rect 429 622 469 624
rect -113 614 -93 620
rect 429 618 465 622
rect 429 617 469 618
rect 429 614 469 615
rect -113 611 -93 612
rect -109 607 -93 611
rect 433 610 469 614
rect 449 598 469 599
rect 54 594 68 598
rect 72 594 74 598
rect 54 592 74 594
rect 449 594 465 598
rect 449 593 469 594
rect 54 589 74 590
rect 54 585 70 589
rect 449 589 469 591
rect 449 585 465 589
rect -113 581 -97 585
rect -113 580 -93 581
rect 54 584 74 585
rect -113 577 -93 578
rect -109 573 -93 577
rect 38 577 74 581
rect 34 576 74 577
rect 34 573 74 574
rect 34 569 70 573
rect 34 568 74 569
rect 34 565 74 566
rect -113 557 -97 561
rect -113 556 -93 557
rect 38 561 74 565
rect 34 560 74 561
rect 34 556 74 558
rect -113 553 -93 554
rect -109 549 -93 553
rect 34 552 70 556
rect 34 551 74 552
rect 34 548 74 549
rect -113 541 -97 545
rect -113 540 -93 541
rect 38 544 74 548
rect -113 537 -93 538
rect -109 533 -93 537
rect 298 537 312 541
rect 316 537 318 541
rect 298 536 318 537
rect 298 533 318 534
rect 54 532 74 533
rect -113 525 -97 529
rect 54 528 70 532
rect -113 524 -93 525
rect 54 527 74 528
rect 302 529 318 533
rect 585 528 601 532
rect 585 527 605 528
rect 54 523 74 525
rect -113 516 -93 522
rect 54 519 70 523
rect 585 524 605 525
rect 589 520 605 524
rect -113 513 -93 514
rect -109 509 -93 513
rect 281 512 316 517
rect 276 511 316 512
rect 276 508 316 509
rect 280 504 316 508
rect 276 503 316 504
rect 585 504 601 508
rect 585 503 605 504
rect 276 500 316 501
rect 276 496 312 500
rect 585 500 605 501
rect 589 496 605 500
rect 280 488 316 492
rect -113 483 -97 487
rect -113 482 -93 483
rect 276 487 316 488
rect 585 488 601 492
rect 276 483 316 485
rect -113 479 -93 480
rect -109 475 -93 479
rect 21 478 35 482
rect 39 478 41 482
rect 21 477 41 478
rect 276 479 312 483
rect 21 474 41 475
rect 25 470 41 474
rect 276 477 316 479
rect 585 487 605 488
rect 585 484 605 485
rect 589 480 605 484
rect 276 474 316 475
rect 281 469 316 474
rect -113 459 -97 463
rect -113 458 -93 459
rect 276 467 316 469
rect 585 472 601 476
rect 585 471 605 472
rect 276 464 316 465
rect 280 460 316 464
rect 585 463 605 469
rect 585 460 605 461
rect -113 455 -93 456
rect -109 451 -93 455
rect 24 453 40 457
rect 20 452 40 453
rect 589 456 605 460
rect 20 447 40 450
rect -113 443 -97 447
rect -113 442 -93 443
rect 20 443 35 447
rect 39 443 40 447
rect -113 439 -93 440
rect -109 435 -93 439
rect 20 440 40 443
rect 449 447 463 451
rect 467 447 469 451
rect 449 445 469 447
rect 449 442 469 443
rect 449 438 465 442
rect 20 437 40 438
rect 24 433 40 437
rect 449 437 469 438
rect -113 427 -97 431
rect 433 430 469 434
rect -113 426 -93 427
rect 429 429 469 430
rect 429 426 469 427
rect -113 418 -93 424
rect 429 422 465 426
rect 429 421 469 422
rect 429 418 469 419
rect -113 415 -93 416
rect -109 411 -93 415
rect 433 414 469 418
rect 429 413 469 414
rect 429 409 469 411
rect 429 405 465 409
rect 429 404 469 405
rect 429 401 469 402
rect 54 396 68 400
rect 72 396 74 400
rect 54 394 74 396
rect 433 397 469 401
rect 54 391 74 392
rect -113 384 -97 388
rect -113 383 -93 384
rect 54 387 70 391
rect 54 386 74 387
rect 449 385 469 386
rect -113 380 -93 381
rect -109 376 -93 380
rect 38 379 74 383
rect 34 378 74 379
rect 449 381 465 385
rect 449 380 469 381
rect 449 376 469 378
rect 34 375 74 376
rect 34 371 70 375
rect -113 360 -97 364
rect -113 359 -93 360
rect 34 370 74 371
rect 449 372 465 376
rect 585 374 601 378
rect 585 373 605 374
rect 585 370 605 371
rect 34 367 74 368
rect 38 363 74 367
rect 34 362 74 363
rect 589 366 605 370
rect 34 358 74 360
rect -113 356 -93 357
rect -109 352 -93 356
rect 34 354 70 358
rect 34 353 74 354
rect 34 350 74 351
rect -113 344 -97 348
rect -113 343 -93 344
rect 38 346 74 350
rect 585 350 601 354
rect 585 349 605 350
rect 585 346 605 347
rect -113 340 -93 341
rect -109 336 -93 340
rect 589 342 605 346
rect 54 334 74 335
rect -113 328 -97 332
rect 54 330 70 334
rect -113 327 -93 328
rect 54 329 74 330
rect 298 332 312 336
rect 316 332 318 336
rect 298 331 318 332
rect 585 334 601 338
rect 585 333 605 334
rect 585 330 605 331
rect 298 328 318 329
rect 54 325 74 327
rect -113 319 -93 325
rect 54 321 70 325
rect 302 324 318 328
rect 589 326 605 330
rect 585 318 601 322
rect -113 316 -93 317
rect -109 312 -93 316
rect 585 317 605 318
rect 279 303 315 307
rect 279 302 319 303
rect 585 309 605 315
rect 585 306 605 307
rect 589 302 605 306
rect 279 298 319 300
rect 279 294 315 298
rect -113 286 -97 290
rect -113 285 -93 286
rect 279 292 319 294
rect 449 293 463 297
rect 467 293 469 297
rect 279 288 319 290
rect -113 282 -93 283
rect -109 278 -93 282
rect 21 281 35 285
rect 39 281 41 285
rect 21 280 41 281
rect 283 284 319 288
rect 279 282 319 284
rect 449 291 469 293
rect 449 288 469 289
rect 449 284 465 288
rect 449 283 469 284
rect 279 279 319 280
rect 21 277 41 278
rect 25 273 41 277
rect 279 275 315 279
rect 433 276 469 280
rect 429 275 469 276
rect 429 272 469 273
rect -113 262 -97 266
rect -113 261 -93 262
rect 429 268 465 272
rect 429 267 469 268
rect 585 266 601 270
rect 585 265 605 266
rect 429 264 469 265
rect 433 260 469 264
rect -113 258 -93 259
rect -109 254 -93 258
rect 24 256 40 260
rect 20 255 40 256
rect 429 259 469 260
rect 585 262 605 263
rect 589 258 605 262
rect 429 255 469 257
rect 20 250 40 253
rect -113 246 -97 250
rect -113 245 -93 246
rect 20 246 35 250
rect 39 246 40 250
rect -113 242 -93 243
rect -109 238 -93 242
rect 20 243 40 246
rect 429 251 465 255
rect 429 250 469 251
rect 429 247 469 248
rect 433 243 469 247
rect 585 242 601 246
rect 585 241 605 242
rect 20 240 40 241
rect 24 236 40 240
rect 585 238 605 239
rect 589 234 605 238
rect -113 230 -97 234
rect 449 231 469 232
rect -113 229 -93 230
rect 449 227 465 231
rect -113 221 -93 227
rect 449 226 469 227
rect 585 226 601 230
rect 449 222 469 224
rect -113 218 -93 219
rect -109 214 -93 218
rect 449 218 465 222
rect 585 225 605 226
rect 585 222 605 223
rect 589 218 605 222
rect 585 210 601 214
rect 585 209 605 210
rect 585 201 605 207
rect 585 198 605 199
rect 54 193 68 197
rect 72 193 74 197
rect -113 189 -97 193
rect -113 188 -93 189
rect 54 191 74 193
rect 589 194 605 198
rect 54 188 74 189
rect -113 185 -93 186
rect -109 181 -93 185
rect 54 184 70 188
rect 54 183 74 184
rect 38 176 74 180
rect -113 165 -97 169
rect -113 164 -93 165
rect 34 175 74 176
rect 34 172 74 173
rect 34 168 70 172
rect 34 167 74 168
rect 34 164 74 165
rect -113 161 -93 162
rect -109 157 -93 161
rect 38 160 74 164
rect 34 159 74 160
rect 34 155 74 157
rect -113 149 -97 153
rect -113 148 -93 149
rect 34 151 70 155
rect -113 145 -93 146
rect -109 141 -93 145
rect 34 150 74 151
rect 34 147 74 148
rect 38 143 74 147
rect -113 133 -97 137
rect -113 132 -93 133
rect 54 131 74 132
rect -113 124 -93 130
rect 54 127 70 131
rect 54 126 74 127
rect 54 122 74 124
rect -113 121 -93 122
rect -109 117 -93 121
rect 54 118 70 122
rect -113 89 -97 93
rect -113 88 -93 89
rect -113 85 -93 86
rect -109 81 -93 85
rect -113 65 -97 69
rect -113 64 -93 65
rect 21 66 35 70
rect 39 66 41 70
rect 21 65 41 66
rect 21 62 41 63
rect -113 61 -93 62
rect -109 57 -93 61
rect 25 58 41 62
rect -113 49 -97 53
rect -113 48 -93 49
rect -113 45 -93 46
rect -109 41 -93 45
rect 24 41 40 45
rect 20 40 40 41
rect -113 33 -97 37
rect 20 35 40 38
rect -113 32 -93 33
rect 20 31 35 35
rect 39 31 40 35
rect -113 24 -93 30
rect 20 28 40 31
rect 20 25 40 26
rect -113 21 -93 22
rect -109 17 -93 21
rect 24 21 40 25
<< ndcontact >>
rect 95 987 99 991
rect 468 990 472 994
rect 474 982 478 986
rect 99 978 103 982
rect -75 974 -71 978
rect 468 974 472 978
rect -69 966 -65 970
rect 91 970 95 974
rect 331 968 335 972
rect -75 958 -71 962
rect 335 960 339 964
rect 474 958 478 962
rect 107 954 111 958
rect -69 942 -65 946
rect 474 950 478 954
rect -69 934 -65 938
rect 91 937 95 941
rect 328 942 332 946
rect 344 933 348 937
rect 468 934 472 938
rect 623 935 627 939
rect -75 918 -71 922
rect 93 921 97 925
rect 344 924 348 928
rect 468 926 472 930
rect 629 927 633 931
rect -75 910 -71 914
rect 99 912 103 916
rect 328 916 332 920
rect 474 918 478 922
rect 623 919 627 923
rect -69 902 -65 906
rect 344 907 348 911
rect 629 903 633 907
rect 328 897 332 901
rect 629 895 633 899
rect 344 887 348 891
rect -75 877 -71 881
rect 344 878 348 882
rect 623 879 627 883
rect -69 869 -65 873
rect 55 872 59 876
rect -75 861 -71 865
rect 59 864 63 868
rect 328 870 332 874
rect 623 871 627 875
rect 344 861 348 865
rect 629 863 633 867
rect -69 845 -65 849
rect 52 847 56 851
rect 490 854 494 858
rect -69 837 -65 841
rect 344 842 348 846
rect 494 845 498 849
rect 486 837 490 841
rect 58 827 62 831
rect -75 821 -71 825
rect 502 821 506 825
rect -75 813 -71 817
rect -69 805 -65 809
rect 486 804 490 808
rect 95 792 99 796
rect 99 783 103 787
rect 488 788 492 792
rect -75 778 -71 782
rect 494 779 498 783
rect -69 770 -65 774
rect 91 775 95 779
rect -75 762 -71 766
rect 107 759 111 763
rect 331 758 335 762
rect -69 746 -65 750
rect 335 750 339 754
rect 91 742 95 746
rect -69 738 -65 742
rect 623 741 627 745
rect -75 722 -71 726
rect 93 726 97 730
rect 328 732 332 736
rect 629 733 633 737
rect -75 714 -71 718
rect 99 717 103 721
rect 344 723 348 727
rect 623 725 627 729
rect -69 706 -65 710
rect 629 709 633 713
rect 328 704 332 708
rect 328 696 332 700
rect 629 701 633 705
rect -75 679 -71 683
rect 328 687 332 691
rect 623 685 627 689
rect 344 678 348 682
rect -69 671 -65 675
rect 55 672 59 676
rect -75 663 -71 667
rect 59 664 63 668
rect 328 670 332 674
rect 623 677 627 681
rect 629 669 633 673
rect 328 661 332 665
rect 344 652 348 656
rect 490 660 494 664
rect 494 651 498 655
rect -69 647 -65 651
rect 52 647 56 651
rect -69 639 -65 643
rect 486 643 490 647
rect 58 627 62 631
rect -75 623 -71 627
rect 502 627 506 631
rect -75 615 -71 619
rect -69 607 -65 611
rect 486 610 490 614
rect 95 594 99 598
rect 488 594 492 598
rect 99 585 103 589
rect 494 585 498 589
rect -75 581 -71 585
rect -69 573 -65 577
rect 91 577 95 581
rect -75 565 -71 569
rect 107 561 111 565
rect -69 549 -65 553
rect -69 541 -65 545
rect 91 544 95 548
rect 332 537 336 541
rect -75 525 -71 529
rect 93 528 97 532
rect 336 529 340 533
rect 623 528 627 532
rect -75 517 -71 521
rect 99 519 103 523
rect 629 520 633 524
rect -69 509 -65 513
rect 330 512 334 516
rect 623 512 627 516
rect 346 504 350 508
rect 346 496 350 500
rect 629 496 633 500
rect -75 483 -71 487
rect 346 488 350 492
rect -69 475 -65 479
rect 55 478 59 482
rect -75 467 -71 471
rect 629 488 633 492
rect 330 479 334 483
rect 59 470 63 474
rect 330 469 334 473
rect 623 472 627 476
rect 346 460 350 464
rect 623 464 627 468
rect -69 451 -65 455
rect 52 453 56 457
rect 629 456 633 460
rect -69 443 -65 447
rect 490 447 494 451
rect 494 438 498 442
rect 58 433 62 437
rect -75 427 -71 431
rect 486 430 490 434
rect -75 419 -71 423
rect -69 411 -65 415
rect 502 414 506 418
rect 95 396 99 400
rect 486 397 490 401
rect -75 384 -71 388
rect 99 387 103 391
rect -69 376 -65 380
rect 91 379 95 383
rect 488 381 492 385
rect -75 368 -71 372
rect 494 372 498 376
rect 623 374 627 378
rect 107 363 111 367
rect 629 366 633 370
rect -69 352 -65 356
rect 623 358 627 362
rect -69 344 -65 348
rect 91 346 95 350
rect 629 342 633 346
rect -75 328 -71 332
rect 93 330 97 334
rect 332 332 336 336
rect 629 334 633 338
rect -75 320 -71 324
rect 99 321 103 325
rect 336 324 340 328
rect 623 318 627 322
rect -69 312 -65 316
rect 349 303 353 307
rect 623 310 627 314
rect 629 302 633 306
rect -75 286 -71 290
rect 333 294 337 298
rect -69 278 -65 282
rect 55 281 59 285
rect 490 293 494 297
rect 494 284 498 288
rect -75 270 -71 274
rect 59 273 63 277
rect 349 275 353 279
rect 486 276 490 280
rect 623 266 627 270
rect -69 254 -65 258
rect 52 256 56 260
rect 502 260 506 264
rect 629 258 633 262
rect -69 246 -65 250
rect 623 250 627 254
rect 486 243 490 247
rect 58 236 62 240
rect 629 234 633 238
rect -75 230 -71 234
rect -75 222 -71 226
rect 488 227 492 231
rect 629 226 633 230
rect 494 218 498 222
rect -69 214 -65 218
rect 623 210 627 214
rect 623 202 627 206
rect -75 189 -71 193
rect 95 193 99 197
rect 629 194 633 198
rect -69 181 -65 185
rect 99 184 103 188
rect -75 173 -71 177
rect 91 176 95 180
rect -69 157 -65 161
rect 107 160 111 164
rect -69 149 -65 153
rect 91 143 95 147
rect -75 133 -71 137
rect -75 125 -71 129
rect 93 127 97 131
rect -69 117 -65 121
rect 99 118 103 122
rect -75 89 -71 93
rect -69 81 -65 85
rect -75 73 -71 77
rect 55 66 59 70
rect -69 57 -65 61
rect 59 58 63 62
rect -69 49 -65 53
rect 52 41 56 45
rect -75 33 -71 37
rect -75 25 -71 29
rect 58 21 62 25
rect -69 17 -65 21
<< pdcontact >>
rect 68 987 72 991
rect 446 990 450 994
rect 70 978 74 982
rect 430 982 434 986
rect -97 974 -93 978
rect -113 966 -109 970
rect 34 970 38 974
rect 311 968 315 972
rect 70 962 74 966
rect 446 966 450 970
rect 297 960 301 964
rect -97 950 -93 954
rect 34 954 38 958
rect 430 958 434 962
rect 128 954 132 958
rect -113 942 -109 946
rect 70 945 74 949
rect 446 950 450 954
rect 310 942 314 946
rect -97 934 -93 938
rect 34 937 38 941
rect 430 942 434 946
rect -113 926 -109 930
rect 274 933 278 937
rect 446 934 450 938
rect 601 935 605 939
rect -97 918 -93 922
rect 70 921 74 925
rect 310 924 314 928
rect 585 927 589 931
rect 70 912 74 916
rect 274 916 278 920
rect 430 918 434 922
rect 274 907 278 911
rect -113 902 -109 906
rect 601 911 605 915
rect 585 903 589 907
rect 310 897 314 901
rect 601 895 605 899
rect 274 887 278 891
rect 585 887 589 891
rect -97 877 -93 881
rect 310 878 314 882
rect 601 879 605 883
rect -113 869 -109 873
rect 35 872 39 876
rect 274 870 278 874
rect 21 864 25 868
rect 274 861 278 865
rect -97 853 -93 857
rect 585 863 589 867
rect 310 851 314 855
rect -113 845 -109 849
rect 20 847 24 851
rect 463 854 467 858
rect -97 837 -93 841
rect 35 837 39 841
rect -113 829 -109 833
rect 274 842 278 846
rect 465 845 469 849
rect 429 837 433 841
rect 20 827 24 831
rect 465 829 469 833
rect -97 821 -93 825
rect 429 821 433 825
rect 523 821 527 825
rect 465 812 469 816
rect -113 805 -109 809
rect 429 804 433 808
rect 68 792 72 796
rect 465 788 469 792
rect 70 783 74 787
rect -97 778 -93 782
rect 465 779 469 783
rect 34 775 38 779
rect -113 770 -109 774
rect 70 767 74 771
rect -97 754 -93 758
rect 34 759 38 763
rect 128 759 132 763
rect 311 758 315 762
rect -113 746 -109 750
rect 70 750 74 754
rect 297 750 301 754
rect 34 742 38 746
rect -97 738 -93 742
rect 601 741 605 745
rect -113 730 -109 734
rect 274 732 278 736
rect 70 726 74 730
rect -97 722 -93 726
rect 585 733 589 737
rect 274 723 278 727
rect 70 717 74 721
rect 310 713 314 717
rect -113 706 -109 710
rect 601 717 605 721
rect 585 709 589 713
rect 274 704 278 708
rect 601 701 605 705
rect 310 696 314 700
rect 585 693 589 697
rect 274 687 278 691
rect -97 679 -93 683
rect 601 685 605 689
rect 274 678 278 682
rect -113 671 -109 675
rect 35 672 39 676
rect 310 670 314 674
rect 21 664 25 668
rect 585 669 589 673
rect -97 655 -93 659
rect 274 661 278 665
rect 463 660 467 664
rect 274 652 278 656
rect -113 647 -109 651
rect 465 651 469 655
rect 20 647 24 651
rect -97 639 -93 643
rect -113 631 -109 635
rect 35 637 39 641
rect 429 643 433 647
rect 465 635 469 639
rect 20 627 24 631
rect 429 627 433 631
rect -97 623 -93 627
rect 523 627 527 631
rect 465 618 469 622
rect -113 607 -109 611
rect 429 610 433 614
rect 68 594 72 598
rect 465 594 469 598
rect 70 585 74 589
rect 465 585 469 589
rect -97 581 -93 585
rect -113 573 -109 577
rect 34 577 38 581
rect 70 569 74 573
rect -97 557 -93 561
rect 34 561 38 565
rect 128 561 132 565
rect -113 549 -109 553
rect 70 552 74 556
rect -97 541 -93 545
rect 34 544 38 548
rect -113 533 -109 537
rect 312 537 316 541
rect -97 525 -93 529
rect 70 528 74 532
rect 298 529 302 533
rect 601 528 605 532
rect 70 519 74 523
rect 585 520 589 524
rect -113 509 -109 513
rect 276 504 280 508
rect 601 504 605 508
rect 312 496 316 500
rect 585 496 589 500
rect 276 488 280 492
rect -97 483 -93 487
rect 601 488 605 492
rect -113 475 -109 479
rect 35 478 39 482
rect 312 479 316 483
rect 21 470 25 474
rect 585 480 589 484
rect -97 459 -93 463
rect 601 472 605 476
rect 276 460 280 464
rect -113 451 -109 455
rect 20 453 24 457
rect 585 456 589 460
rect -97 443 -93 447
rect 35 443 39 447
rect -113 435 -109 439
rect 463 447 467 451
rect 465 438 469 442
rect 20 433 24 437
rect -97 427 -93 431
rect 429 430 433 434
rect 465 422 469 426
rect -113 411 -109 415
rect 429 414 433 418
rect 523 414 527 418
rect 465 405 469 409
rect 68 396 72 400
rect 429 397 433 401
rect -97 384 -93 388
rect 70 387 74 391
rect -113 376 -109 380
rect 34 379 38 383
rect 465 381 469 385
rect 70 371 74 375
rect -97 360 -93 364
rect 465 372 469 376
rect 601 374 605 378
rect 34 363 38 367
rect 128 363 132 367
rect 585 366 589 370
rect -113 352 -109 356
rect 70 354 74 358
rect -97 344 -93 348
rect 34 346 38 350
rect 601 350 605 354
rect -113 336 -109 340
rect 585 342 589 346
rect -97 328 -93 332
rect 70 330 74 334
rect 312 332 316 336
rect 601 334 605 338
rect 70 321 74 325
rect 298 324 302 328
rect 585 326 589 330
rect 601 318 605 322
rect -113 312 -109 316
rect 315 303 319 307
rect 585 302 589 306
rect 315 294 319 298
rect -97 286 -93 290
rect 463 293 467 297
rect -113 278 -109 282
rect 35 281 39 285
rect 279 284 283 288
rect 465 284 469 288
rect 21 273 25 277
rect 315 275 319 279
rect 429 276 433 280
rect -97 262 -93 266
rect 465 268 469 272
rect 601 266 605 270
rect 429 260 433 264
rect -113 254 -109 258
rect 20 256 24 260
rect 523 260 527 264
rect 585 258 589 262
rect -97 246 -93 250
rect 35 246 39 250
rect -113 238 -109 242
rect 465 251 469 255
rect 429 243 433 247
rect 601 242 605 246
rect 20 236 24 240
rect 585 234 589 238
rect -97 230 -93 234
rect 465 227 469 231
rect 601 226 605 230
rect -113 214 -109 218
rect 465 218 469 222
rect 585 218 589 222
rect 601 210 605 214
rect 68 193 72 197
rect -97 189 -93 193
rect 585 194 589 198
rect -113 181 -109 185
rect 70 184 74 188
rect 34 176 38 180
rect -97 165 -93 169
rect 70 168 74 172
rect -113 157 -109 161
rect 34 160 38 164
rect 128 160 132 164
rect -97 149 -93 153
rect 70 151 74 155
rect -113 141 -109 145
rect 34 143 38 147
rect -97 133 -93 137
rect 70 127 74 131
rect -113 117 -109 121
rect 70 118 74 122
rect -97 89 -93 93
rect -113 81 -109 85
rect -97 65 -93 69
rect 35 66 39 70
rect -113 57 -109 61
rect 21 58 25 62
rect -97 49 -93 53
rect -113 41 -109 45
rect 20 41 24 45
rect -97 33 -93 37
rect 35 31 39 35
rect -113 17 -109 21
rect 20 21 24 25
<< psubstratepcontact >>
rect 343 960 347 964
rect 115 954 119 958
rect 483 918 487 922
rect -60 902 -56 906
rect 67 864 71 868
rect 638 863 642 867
rect 352 842 356 846
rect 66 827 70 831
rect 510 821 514 825
rect -60 805 -56 809
rect 115 759 119 763
rect 343 750 347 754
rect -60 706 -56 710
rect 67 664 71 668
rect 638 669 642 673
rect 352 660 356 664
rect 66 627 70 631
rect 510 627 514 631
rect -60 607 -56 611
rect 115 561 119 565
rect 344 529 348 533
rect -60 509 -56 513
rect 67 470 71 474
rect 354 464 358 468
rect 638 456 642 460
rect 66 433 70 437
rect -60 411 -56 415
rect 510 414 514 418
rect 115 363 119 367
rect 344 324 348 328
rect -60 312 -56 316
rect 638 302 642 306
rect 357 284 361 288
rect 67 273 71 277
rect 510 260 514 264
rect 66 236 70 240
rect -60 214 -56 218
rect 638 194 642 198
rect 115 160 119 164
rect -60 117 -56 121
rect 67 58 71 62
rect 66 21 70 25
rect -60 17 -56 21
<< nsubstratencontact >>
rect 430 974 434 978
rect -113 958 -109 962
rect 289 960 293 964
rect 585 919 589 923
rect 70 902 74 906
rect -113 861 -109 865
rect 13 864 17 868
rect 12 837 16 841
rect 266 842 270 846
rect -113 762 -109 766
rect 465 769 469 773
rect 289 750 293 754
rect 585 725 589 729
rect 70 707 74 711
rect -113 663 -109 667
rect 13 664 17 668
rect 266 652 270 656
rect 12 637 16 641
rect 465 575 469 579
rect -113 565 -109 569
rect 290 529 294 533
rect 70 509 74 513
rect 585 512 589 516
rect -113 467 -109 471
rect 13 470 17 474
rect 268 460 272 464
rect 12 443 16 447
rect -113 368 -109 372
rect 465 362 469 366
rect 585 358 589 362
rect 290 324 294 328
rect 70 311 74 315
rect 271 284 275 288
rect -113 270 -109 274
rect 13 273 17 277
rect 12 246 16 250
rect 585 250 589 254
rect 465 208 469 212
rect -113 173 -109 177
rect 70 108 74 112
rect -113 73 -109 77
rect 13 58 17 62
rect 12 31 16 35
<< polysilicon >>
rect 427 987 430 989
rect 450 987 468 989
rect 478 987 481 989
rect 53 983 54 985
rect 74 983 93 985
rect 103 983 106 985
rect -116 971 -113 973
rect -93 971 -75 973
rect -65 971 -62 973
rect 6 967 34 969
rect 74 967 91 969
rect 111 967 114 969
rect 465 971 468 973
rect 478 971 490 973
rect 294 965 297 967
rect 317 965 329 967
rect 339 965 342 967
rect 22 959 34 961
rect 74 959 91 961
rect 111 959 114 961
rect 427 963 430 965
rect 450 963 468 965
rect 478 963 481 965
rect -78 955 -75 957
rect -65 955 -53 957
rect 5 951 34 953
rect 74 951 91 953
rect 111 951 114 953
rect -116 947 -113 949
rect -93 947 -75 949
rect -65 947 -62 949
rect 419 947 430 949
rect 450 947 468 949
rect 478 947 490 949
rect 6 942 34 944
rect 74 942 91 944
rect 111 942 114 944
rect 263 939 274 941
rect 314 939 328 941
rect 348 939 351 941
rect -124 931 -113 933
rect -93 931 -75 933
rect -65 931 -53 933
rect 458 939 468 941
rect 478 939 481 941
rect 263 929 274 931
rect 314 929 328 931
rect 348 929 351 931
rect 419 931 430 933
rect 450 931 453 933
rect 582 932 585 934
rect 605 932 623 934
rect 633 932 636 934
rect -85 923 -75 925
rect -65 923 -62 925
rect 419 923 430 925
rect 450 923 468 925
rect 478 923 481 925
rect 53 918 54 920
rect 74 918 93 920
rect 103 918 106 920
rect -124 915 -113 917
rect -93 915 -90 917
rect 620 916 623 918
rect 633 916 645 918
rect 263 913 274 915
rect 314 913 328 915
rect 348 913 351 915
rect -124 907 -113 909
rect -93 907 -75 909
rect -65 907 -62 909
rect 582 908 585 910
rect 605 908 623 910
rect 633 908 636 910
rect 263 903 274 905
rect 314 903 328 905
rect 348 903 351 905
rect 263 893 274 895
rect 314 893 328 895
rect 348 893 351 895
rect 574 892 585 894
rect 605 892 623 894
rect 633 892 645 894
rect 263 883 274 885
rect 314 883 328 885
rect 348 883 351 885
rect 613 884 623 886
rect 633 884 636 886
rect -116 874 -113 876
rect -93 874 -75 876
rect -65 874 -62 876
rect 574 876 585 878
rect 605 876 608 878
rect 18 869 21 871
rect 41 869 53 871
rect 63 869 66 871
rect 263 867 274 869
rect 314 867 328 869
rect 348 867 351 869
rect 574 868 585 870
rect 605 868 623 870
rect 633 868 636 870
rect -78 858 -75 860
rect -65 858 -53 860
rect 263 857 274 859
rect 314 857 328 859
rect 348 857 351 859
rect -116 850 -113 852
rect -93 850 -75 852
rect -65 850 -62 852
rect 448 850 449 852
rect 469 850 488 852
rect 498 850 501 852
rect 263 847 274 849
rect 314 847 328 849
rect 348 847 351 849
rect 9 844 20 846
rect 40 844 52 846
rect 62 844 65 846
rect -124 834 -113 836
rect -93 834 -75 836
rect -65 834 -53 836
rect 9 832 20 834
rect 40 832 52 834
rect 62 832 65 834
rect 401 834 429 836
rect 469 834 486 836
rect 506 834 509 836
rect -85 826 -75 828
rect -65 826 -62 828
rect 417 826 429 828
rect 469 826 486 828
rect 506 826 509 828
rect -124 818 -113 820
rect -93 818 -90 820
rect 400 818 429 820
rect 469 818 486 820
rect 506 818 509 820
rect -124 810 -113 812
rect -93 810 -75 812
rect -65 810 -62 812
rect 401 809 429 811
rect 469 809 486 811
rect 506 809 509 811
rect 53 788 54 790
rect 74 788 93 790
rect 103 788 106 790
rect 448 785 449 787
rect 469 785 488 787
rect 498 785 501 787
rect -116 775 -113 777
rect -93 775 -75 777
rect -65 775 -62 777
rect 6 772 34 774
rect 74 772 91 774
rect 111 772 114 774
rect 22 764 34 766
rect 74 764 91 766
rect 111 764 114 766
rect -78 759 -75 761
rect -65 759 -53 761
rect 5 756 34 758
rect 74 756 91 758
rect 111 756 114 758
rect -116 751 -113 753
rect -93 751 -75 753
rect -65 751 -62 753
rect 294 755 297 757
rect 317 755 329 757
rect 339 755 342 757
rect 6 747 34 749
rect 74 747 91 749
rect 111 747 114 749
rect 582 738 585 740
rect 605 738 623 740
rect 633 738 636 740
rect -124 735 -113 737
rect -93 735 -75 737
rect -65 735 -53 737
rect -85 727 -75 729
rect -65 727 -62 729
rect 263 729 274 731
rect 314 729 328 731
rect 348 729 351 731
rect 53 723 54 725
rect 74 723 93 725
rect 103 723 106 725
rect -124 719 -113 721
rect -93 719 -90 721
rect 620 722 623 724
rect 633 722 645 724
rect 263 719 274 721
rect 314 719 328 721
rect 348 719 351 721
rect -124 711 -113 713
rect -93 711 -75 713
rect -65 711 -62 713
rect 582 714 585 716
rect 605 714 623 716
rect 633 714 636 716
rect 263 709 274 711
rect 314 709 328 711
rect 348 709 351 711
rect 574 698 585 700
rect 605 698 623 700
rect 633 698 645 700
rect 263 693 274 695
rect 314 693 328 695
rect 348 693 351 695
rect 613 690 623 692
rect 633 690 636 692
rect 263 683 274 685
rect 314 683 328 685
rect 348 683 351 685
rect 574 682 585 684
rect 605 682 608 684
rect -116 676 -113 678
rect -93 676 -75 678
rect -65 676 -62 678
rect 18 669 21 671
rect 41 669 53 671
rect 63 669 66 671
rect 574 674 585 676
rect 605 674 623 676
rect 633 674 636 676
rect 263 667 274 669
rect 314 667 328 669
rect 348 667 351 669
rect -78 660 -75 662
rect -65 660 -53 662
rect 263 657 274 659
rect 314 657 328 659
rect 348 657 351 659
rect -116 652 -113 654
rect -93 652 -75 654
rect -65 652 -62 654
rect 448 656 449 658
rect 469 656 488 658
rect 498 656 501 658
rect 9 644 20 646
rect 40 644 52 646
rect 62 644 65 646
rect -124 636 -113 638
rect -93 636 -75 638
rect -65 636 -53 638
rect 401 640 429 642
rect 469 640 486 642
rect 506 640 509 642
rect 9 632 20 634
rect 40 632 52 634
rect 62 632 65 634
rect -85 628 -75 630
rect -65 628 -62 630
rect 417 632 429 634
rect 469 632 486 634
rect 506 632 509 634
rect 400 624 429 626
rect 469 624 486 626
rect 506 624 509 626
rect -124 620 -113 622
rect -93 620 -90 622
rect 401 615 429 617
rect 469 615 486 617
rect 506 615 509 617
rect -124 612 -113 614
rect -93 612 -75 614
rect -65 612 -62 614
rect 53 590 54 592
rect 74 590 93 592
rect 103 590 106 592
rect 448 591 449 593
rect 469 591 488 593
rect 498 591 501 593
rect -116 578 -113 580
rect -93 578 -75 580
rect -65 578 -62 580
rect 6 574 34 576
rect 74 574 91 576
rect 111 574 114 576
rect 22 566 34 568
rect 74 566 91 568
rect 111 566 114 568
rect -78 562 -75 564
rect -65 562 -53 564
rect 5 558 34 560
rect 74 558 91 560
rect 111 558 114 560
rect -116 554 -113 556
rect -93 554 -75 556
rect -65 554 -62 556
rect 6 549 34 551
rect 74 549 91 551
rect 111 549 114 551
rect -124 538 -113 540
rect -93 538 -75 540
rect -65 538 -53 540
rect 295 534 298 536
rect 318 534 330 536
rect 340 534 343 536
rect -85 530 -75 532
rect -65 530 -62 532
rect 53 525 54 527
rect 74 525 93 527
rect 103 525 106 527
rect 582 525 585 527
rect 605 525 623 527
rect 633 525 636 527
rect -124 522 -113 524
rect -93 522 -90 524
rect -124 514 -113 516
rect -93 514 -75 516
rect -65 514 -62 516
rect 264 509 276 511
rect 316 509 330 511
rect 350 509 353 511
rect 620 509 623 511
rect 633 509 645 511
rect 264 501 276 503
rect 316 501 330 503
rect 350 501 353 503
rect 582 501 585 503
rect 605 501 623 503
rect 633 501 636 503
rect 264 485 276 487
rect 316 485 330 487
rect 350 485 353 487
rect -116 480 -113 482
rect -93 480 -75 482
rect -65 480 -62 482
rect 18 475 21 477
rect 41 475 53 477
rect 63 475 66 477
rect 574 485 585 487
rect 605 485 623 487
rect 633 485 645 487
rect 264 475 276 477
rect 316 475 330 477
rect 350 475 353 477
rect 613 477 623 479
rect 633 477 636 479
rect -78 464 -75 466
rect -65 464 -53 466
rect 574 469 585 471
rect 605 469 608 471
rect 264 465 276 467
rect 316 465 330 467
rect 350 465 353 467
rect 574 461 585 463
rect 605 461 623 463
rect 633 461 636 463
rect -116 456 -113 458
rect -93 456 -75 458
rect -65 456 -62 458
rect 9 450 20 452
rect 40 450 52 452
rect 62 450 65 452
rect -124 440 -113 442
rect -93 440 -75 442
rect -65 440 -53 442
rect 448 443 449 445
rect 469 443 488 445
rect 498 443 501 445
rect 9 438 20 440
rect 40 438 52 440
rect 62 438 65 440
rect -85 432 -75 434
rect -65 432 -62 434
rect 401 427 429 429
rect 469 427 486 429
rect 506 427 509 429
rect -124 424 -113 426
rect -93 424 -90 426
rect 417 419 429 421
rect 469 419 486 421
rect 506 419 509 421
rect -124 416 -113 418
rect -93 416 -75 418
rect -65 416 -62 418
rect 400 411 429 413
rect 469 411 486 413
rect 506 411 509 413
rect 401 402 429 404
rect 469 402 486 404
rect 506 402 509 404
rect 53 392 54 394
rect 74 392 93 394
rect 103 392 106 394
rect -116 381 -113 383
rect -93 381 -75 383
rect -65 381 -62 383
rect 6 376 34 378
rect 74 376 91 378
rect 111 376 114 378
rect 448 378 449 380
rect 469 378 488 380
rect 498 378 501 380
rect -78 365 -75 367
rect -65 365 -53 367
rect 582 371 585 373
rect 605 371 623 373
rect 633 371 636 373
rect 22 368 34 370
rect 74 368 91 370
rect 111 368 114 370
rect 5 360 34 362
rect 74 360 91 362
rect 111 360 114 362
rect -116 357 -113 359
rect -93 357 -75 359
rect -65 357 -62 359
rect 620 355 623 357
rect 633 355 645 357
rect 6 351 34 353
rect 74 351 91 353
rect 111 351 114 353
rect 582 347 585 349
rect 605 347 623 349
rect 633 347 636 349
rect -124 341 -113 343
rect -93 341 -75 343
rect -65 341 -53 343
rect -85 333 -75 335
rect -65 333 -62 335
rect -124 325 -113 327
rect -93 325 -90 327
rect 295 329 298 331
rect 318 329 330 331
rect 340 329 343 331
rect 574 331 585 333
rect 605 331 623 333
rect 633 331 645 333
rect 53 327 54 329
rect 74 327 93 329
rect 103 327 106 329
rect 613 323 623 325
rect 633 323 636 325
rect -124 317 -113 319
rect -93 317 -75 319
rect -65 317 -62 319
rect 574 315 585 317
rect 605 315 608 317
rect 574 307 585 309
rect 605 307 623 309
rect 633 307 636 309
rect 268 300 279 302
rect 319 300 333 302
rect 353 300 356 302
rect 268 290 279 292
rect 319 290 333 292
rect 353 290 356 292
rect -116 283 -113 285
rect -93 283 -75 285
rect -65 283 -62 285
rect 18 278 21 280
rect 41 278 53 280
rect 63 278 66 280
rect 448 289 449 291
rect 469 289 488 291
rect 498 289 501 291
rect 268 280 279 282
rect 319 280 333 282
rect 353 280 356 282
rect 401 273 429 275
rect 469 273 486 275
rect 506 273 509 275
rect -78 267 -75 269
rect -65 267 -53 269
rect 417 265 429 267
rect 469 265 486 267
rect 506 265 509 267
rect -116 259 -113 261
rect -93 259 -75 261
rect -65 259 -62 261
rect 582 263 585 265
rect 605 263 623 265
rect 633 263 636 265
rect 400 257 429 259
rect 469 257 486 259
rect 506 257 509 259
rect 9 253 20 255
rect 40 253 52 255
rect 62 253 65 255
rect -124 243 -113 245
rect -93 243 -75 245
rect -65 243 -53 245
rect 401 248 429 250
rect 469 248 486 250
rect 506 248 509 250
rect 620 247 623 249
rect 633 247 645 249
rect 9 241 20 243
rect 40 241 52 243
rect 62 241 65 243
rect -85 235 -75 237
rect -65 235 -62 237
rect 582 239 585 241
rect 605 239 623 241
rect 633 239 636 241
rect -124 227 -113 229
rect -93 227 -90 229
rect 448 224 449 226
rect 469 224 488 226
rect 498 224 501 226
rect -124 219 -113 221
rect -93 219 -75 221
rect -65 219 -62 221
rect 574 223 585 225
rect 605 223 623 225
rect 633 223 645 225
rect 613 215 623 217
rect 633 215 636 217
rect 574 207 585 209
rect 605 207 608 209
rect 574 199 585 201
rect 605 199 623 201
rect 633 199 636 201
rect 53 189 54 191
rect 74 189 93 191
rect 103 189 106 191
rect -116 186 -113 188
rect -93 186 -75 188
rect -65 186 -62 188
rect -78 170 -75 172
rect -65 170 -53 172
rect 6 173 34 175
rect 74 173 91 175
rect 111 173 114 175
rect 22 165 34 167
rect 74 165 91 167
rect 111 165 114 167
rect -116 162 -113 164
rect -93 162 -75 164
rect -65 162 -62 164
rect 5 157 34 159
rect 74 157 91 159
rect 111 157 114 159
rect -124 146 -113 148
rect -93 146 -75 148
rect -65 146 -53 148
rect 6 148 34 150
rect 74 148 91 150
rect 111 148 114 150
rect -85 138 -75 140
rect -65 138 -62 140
rect -124 130 -113 132
rect -93 130 -90 132
rect -124 122 -113 124
rect -93 122 -75 124
rect -65 122 -62 124
rect 53 124 54 126
rect 74 124 93 126
rect 103 124 106 126
rect -116 86 -113 88
rect -93 86 -75 88
rect -65 86 -62 88
rect -78 70 -75 72
rect -65 70 -53 72
rect -116 62 -113 64
rect -93 62 -75 64
rect -65 62 -62 64
rect 18 63 21 65
rect 41 63 53 65
rect 63 63 66 65
rect -124 46 -113 48
rect -93 46 -75 48
rect -65 46 -53 48
rect -85 38 -75 40
rect -65 38 -62 40
rect 9 38 20 40
rect 40 38 52 40
rect 62 38 65 40
rect -124 30 -113 32
rect -93 30 -90 32
rect 9 26 20 28
rect 40 26 52 28
rect 62 26 65 28
rect -124 22 -113 24
rect -93 22 -75 24
rect -65 22 -62 24
<< polycontact >>
rect 49 982 53 986
rect 459 983 463 987
rect -84 967 -80 971
rect 2 966 6 970
rect 18 958 22 962
rect 490 970 494 974
rect 320 961 324 965
rect -53 954 -49 958
rect 1 950 5 954
rect 460 959 464 963
rect -83 943 -79 947
rect 2 941 6 945
rect 415 946 419 950
rect -128 930 -124 934
rect 259 938 263 942
rect -89 922 -85 926
rect -53 930 -49 934
rect 259 928 263 932
rect 454 938 458 942
rect 490 946 494 950
rect 415 930 419 934
rect -128 914 -124 918
rect 49 917 53 921
rect 415 922 419 926
rect 614 928 618 932
rect -128 906 -124 910
rect 259 912 263 916
rect 259 902 263 906
rect 645 915 649 919
rect 615 904 619 908
rect 259 892 263 896
rect 259 882 263 886
rect 570 891 574 895
rect 609 883 613 887
rect 645 891 649 895
rect -84 870 -80 874
rect 570 875 574 879
rect 44 865 48 869
rect 259 866 263 870
rect 570 867 574 871
rect -53 857 -49 861
rect 259 856 263 860
rect -83 846 -79 850
rect 5 843 9 847
rect 259 846 263 850
rect 444 849 448 853
rect -128 833 -124 837
rect -89 825 -85 829
rect -53 833 -49 837
rect 5 831 9 835
rect 397 833 401 837
rect 413 825 417 829
rect -128 817 -124 821
rect -128 809 -124 813
rect 396 817 400 821
rect 397 808 401 812
rect 49 787 53 791
rect 444 784 448 788
rect -84 771 -80 775
rect 2 771 6 775
rect 18 763 22 767
rect -53 758 -49 762
rect 1 755 5 759
rect -83 747 -79 751
rect 2 746 6 750
rect 320 751 324 755
rect -128 734 -124 738
rect -89 726 -85 730
rect -53 734 -49 738
rect 49 722 53 726
rect 259 728 263 732
rect 614 734 618 738
rect -128 718 -124 722
rect -128 710 -124 714
rect 259 718 263 722
rect 259 708 263 712
rect 645 721 649 725
rect 615 710 619 714
rect 259 692 263 696
rect 570 697 574 701
rect 259 682 263 686
rect 609 689 613 693
rect 645 697 649 701
rect 570 681 574 685
rect -84 672 -80 676
rect 44 665 48 669
rect 259 666 263 670
rect 570 673 574 677
rect -53 659 -49 663
rect 259 656 263 660
rect 444 655 448 659
rect -83 648 -79 652
rect 5 643 9 647
rect -128 635 -124 639
rect -89 627 -85 631
rect -53 635 -49 639
rect 5 631 9 635
rect 397 639 401 643
rect 413 631 417 635
rect 396 623 400 627
rect -128 619 -124 623
rect -128 611 -124 615
rect 397 614 401 618
rect 49 589 53 593
rect 444 590 448 594
rect -84 574 -80 578
rect 2 573 6 577
rect 18 565 22 569
rect -53 561 -49 565
rect 1 557 5 561
rect -83 550 -79 554
rect 2 548 6 552
rect -128 537 -124 541
rect -89 529 -85 533
rect -53 537 -49 541
rect -128 521 -124 525
rect 49 524 53 528
rect 321 530 325 534
rect -128 513 -124 517
rect 614 521 618 525
rect 260 508 264 512
rect 260 500 264 504
rect 645 508 649 512
rect 615 497 619 501
rect 260 484 264 488
rect -84 476 -80 480
rect 44 471 48 475
rect 260 474 264 478
rect 570 484 574 488
rect 609 476 613 480
rect 645 484 649 488
rect -53 463 -49 467
rect 260 464 264 468
rect 570 468 574 472
rect 570 460 574 464
rect -83 452 -79 456
rect 5 449 9 453
rect -128 439 -124 443
rect -89 431 -85 435
rect -53 439 -49 443
rect 5 437 9 441
rect 444 442 448 446
rect -128 423 -124 427
rect 397 426 401 430
rect -128 415 -124 419
rect 413 418 417 422
rect 396 410 400 414
rect 397 401 401 405
rect 49 391 53 395
rect -84 377 -80 381
rect 2 375 6 379
rect 444 377 448 381
rect -53 364 -49 368
rect 18 367 22 371
rect 1 359 5 363
rect 614 367 618 371
rect -83 353 -79 357
rect 2 350 6 354
rect -128 340 -124 344
rect 645 354 649 358
rect -89 332 -85 336
rect -53 340 -49 344
rect 615 343 619 347
rect -128 324 -124 328
rect 49 326 53 330
rect 570 330 574 334
rect -128 316 -124 320
rect 321 325 325 329
rect 609 322 613 326
rect 645 330 649 334
rect 570 314 574 318
rect 264 299 268 303
rect 570 306 574 310
rect 264 289 268 293
rect -84 279 -80 283
rect 264 279 268 283
rect 444 288 448 292
rect 44 274 48 278
rect 397 272 401 276
rect -53 266 -49 270
rect 413 264 417 268
rect -83 255 -79 259
rect 5 252 9 256
rect 396 256 400 260
rect 614 259 618 263
rect -128 242 -124 246
rect -89 234 -85 238
rect -53 242 -49 246
rect 5 240 9 244
rect 397 247 401 251
rect 645 246 649 250
rect 615 235 619 239
rect -128 226 -124 230
rect -128 218 -124 222
rect 444 223 448 227
rect 570 222 574 226
rect 609 214 613 218
rect 645 222 649 226
rect 570 206 574 210
rect 570 198 574 202
rect 49 188 53 192
rect -84 182 -80 186
rect -53 169 -49 173
rect 2 172 6 176
rect 18 164 22 168
rect -83 158 -79 162
rect 1 156 5 160
rect -128 145 -124 149
rect -89 137 -85 141
rect -53 145 -49 149
rect 2 147 6 151
rect -128 129 -124 133
rect -128 121 -124 125
rect 49 123 53 127
rect -84 82 -80 86
rect -53 69 -49 73
rect -83 58 -79 62
rect 44 59 48 63
rect -128 45 -124 49
rect -89 37 -85 41
rect -53 45 -49 49
rect 5 37 9 41
rect -128 29 -124 33
rect -128 21 -124 25
rect 5 25 9 29
<< metal1 >>
rect -121 1030 581 1034
rect -121 970 -117 1030
rect -82 978 -78 986
rect -93 974 -75 978
rect -121 966 -113 970
rect -121 962 -117 966
rect -84 962 -80 967
rect -65 966 -33 970
rect -121 958 -113 962
rect -89 959 -75 962
rect -121 946 -117 958
rect -89 954 -86 959
rect -93 950 -86 954
rect -121 942 -113 946
rect -60 946 -56 966
rect -128 918 -124 930
rect -139 914 -128 918
rect -121 930 -117 942
rect -83 938 -79 943
rect -65 942 -56 946
rect -60 938 -56 942
rect -93 934 -79 938
rect -65 934 -56 938
rect -121 926 -113 930
rect -139 821 -135 914
rect -121 906 -117 926
rect -93 918 -85 922
rect -82 922 -79 934
rect -82 918 -75 922
rect -88 914 -85 918
rect -88 910 -75 914
rect -60 906 -56 934
rect -53 934 -49 954
rect -121 902 -113 906
rect -65 902 -60 906
rect -121 873 -117 902
rect -82 881 -78 886
rect -93 877 -75 881
rect -121 869 -113 873
rect -37 873 -33 966
rect -121 865 -117 869
rect -84 865 -80 870
rect -65 869 -33 873
rect -121 861 -113 865
rect -89 862 -75 865
rect -121 849 -117 861
rect -89 857 -86 862
rect -93 853 -86 857
rect -121 845 -113 849
rect -60 849 -56 869
rect -128 821 -124 833
rect -139 817 -128 821
rect -121 833 -117 845
rect -83 841 -79 846
rect -65 845 -56 849
rect -60 841 -56 845
rect -93 837 -79 841
rect -65 837 -56 841
rect -121 829 -113 833
rect -139 722 -135 817
rect -121 809 -117 829
rect -93 821 -85 825
rect -82 825 -79 837
rect -82 821 -75 825
rect -88 817 -85 821
rect -88 813 -75 817
rect -60 809 -56 837
rect -53 837 -49 857
rect -121 805 -113 809
rect -65 805 -60 809
rect -121 774 -117 805
rect -82 782 -78 786
rect -93 778 -75 782
rect -121 770 -113 774
rect -37 774 -33 869
rect -29 962 -25 986
rect -29 848 -25 957
rect -21 891 -17 941
rect -21 836 -17 886
rect -13 906 -9 1030
rect 2 994 81 998
rect 2 970 6 994
rect 77 991 81 994
rect 72 987 95 991
rect 10 982 49 986
rect 1 954 5 957
rect 10 945 14 982
rect 74 978 77 982
rect 103 978 119 982
rect 26 970 34 974
rect 6 941 14 945
rect 18 933 22 958
rect 26 958 30 970
rect 86 966 90 970
rect 74 962 90 966
rect 26 954 34 958
rect 26 941 30 954
rect 74 945 77 949
rect 86 941 90 962
rect 115 958 119 978
rect 111 954 115 958
rect 119 954 128 958
rect 132 954 156 958
rect 26 937 34 941
rect 86 937 91 941
rect 18 929 89 933
rect 85 925 89 929
rect 74 921 93 925
rect 14 917 49 921
rect 74 912 77 916
rect 115 916 119 954
rect 103 912 119 916
rect 70 906 74 912
rect -13 902 70 906
rect -13 868 -9 902
rect 44 876 48 879
rect 39 872 55 876
rect -13 864 13 868
rect 17 864 21 868
rect 152 868 156 954
rect -121 766 -117 770
rect -84 766 -80 771
rect -65 770 -33 774
rect -121 762 -113 766
rect -89 763 -75 766
rect -121 750 -117 762
rect -89 758 -86 763
rect -93 754 -86 758
rect -121 746 -113 750
rect -60 750 -56 770
rect -128 722 -124 734
rect -139 718 -128 722
rect -121 734 -117 746
rect -83 742 -79 747
rect -65 746 -56 750
rect -60 742 -56 746
rect -93 738 -79 742
rect -65 738 -56 742
rect -121 730 -113 734
rect -139 623 -135 718
rect -121 710 -117 730
rect -93 722 -85 726
rect -82 726 -79 738
rect -82 722 -75 726
rect -88 718 -85 722
rect -88 714 -75 718
rect -60 710 -56 738
rect -53 738 -49 758
rect -121 706 -113 710
rect -65 706 -60 710
rect -121 675 -117 706
rect -82 683 -78 686
rect -93 679 -75 683
rect -121 671 -113 675
rect -37 675 -33 770
rect -121 667 -117 671
rect -84 667 -80 672
rect -65 671 -33 675
rect -121 663 -113 667
rect -89 664 -75 667
rect -121 651 -117 663
rect -89 659 -86 664
rect -93 655 -86 659
rect -121 647 -113 651
rect -60 651 -56 671
rect -128 623 -124 635
rect -139 619 -128 623
rect -121 635 -117 647
rect -83 643 -79 648
rect -65 647 -56 651
rect -60 643 -56 647
rect -93 639 -79 643
rect -65 639 -56 643
rect -121 631 -113 635
rect -139 525 -135 619
rect -121 611 -117 631
rect -93 623 -85 627
rect -82 627 -79 639
rect -82 623 -75 627
rect -88 619 -85 623
rect -88 615 -75 619
rect -60 611 -56 639
rect -53 639 -49 659
rect -121 607 -113 611
rect -65 607 -60 611
rect -121 577 -117 607
rect -82 585 -78 590
rect -93 581 -75 585
rect -121 573 -113 577
rect -37 577 -33 671
rect -29 767 -25 786
rect -29 648 -25 762
rect -21 691 -17 746
rect -21 636 -17 686
rect -13 711 -9 864
rect 12 851 16 864
rect 44 851 48 865
rect 63 864 67 868
rect 71 864 156 868
rect 12 847 20 851
rect 44 847 52 851
rect 4 843 5 847
rect 12 841 16 847
rect 44 841 48 847
rect 39 837 48 841
rect 4 831 5 835
rect 12 831 16 837
rect 152 831 156 864
rect 12 827 20 831
rect 62 827 66 831
rect 70 827 156 831
rect 2 799 81 803
rect 2 775 6 799
rect 77 796 81 799
rect 72 792 95 796
rect 10 787 49 791
rect 1 759 5 762
rect 10 750 14 787
rect 74 783 77 787
rect 103 783 119 787
rect 26 775 34 779
rect 6 746 14 750
rect 18 738 22 763
rect 26 763 30 775
rect 86 771 90 775
rect 74 767 90 771
rect 26 759 34 763
rect 26 746 30 759
rect 74 750 77 754
rect 86 746 90 767
rect 115 763 119 783
rect 152 763 156 827
rect 111 759 115 763
rect 119 759 128 763
rect 132 759 156 763
rect 26 742 34 746
rect 86 742 91 746
rect 18 734 89 738
rect 85 730 89 734
rect 74 726 93 730
rect 14 722 49 726
rect 74 717 77 721
rect 115 721 119 759
rect 103 717 119 721
rect 70 711 74 717
rect -13 707 70 711
rect -13 668 -9 707
rect 44 676 48 679
rect 39 672 55 676
rect -13 664 13 668
rect 17 664 21 668
rect 152 668 156 759
rect -121 569 -117 573
rect -84 569 -80 574
rect -65 573 -33 577
rect -121 565 -113 569
rect -89 566 -75 569
rect -121 553 -117 565
rect -89 561 -86 566
rect -93 557 -86 561
rect -121 549 -113 553
rect -60 553 -56 573
rect -128 525 -124 537
rect -139 521 -128 525
rect -121 537 -117 549
rect -83 545 -79 550
rect -65 549 -56 553
rect -60 545 -56 549
rect -93 541 -79 545
rect -65 541 -56 545
rect -121 533 -113 537
rect -139 427 -135 521
rect -121 513 -117 533
rect -93 525 -85 529
rect -82 529 -79 541
rect -82 525 -75 529
rect -88 521 -85 525
rect -88 517 -75 521
rect -60 513 -56 541
rect -53 541 -49 561
rect -121 509 -113 513
rect -65 509 -60 513
rect -121 479 -117 509
rect -82 487 -78 492
rect -93 483 -75 487
rect -121 475 -113 479
rect -37 479 -33 573
rect -121 471 -117 475
rect -84 471 -80 476
rect -65 475 -33 479
rect -121 467 -113 471
rect -89 468 -75 471
rect -121 455 -117 467
rect -89 463 -86 468
rect -93 459 -86 463
rect -121 451 -113 455
rect -60 455 -56 475
rect -128 427 -124 439
rect -139 423 -128 427
rect -121 439 -117 451
rect -83 447 -79 452
rect -65 451 -56 455
rect -60 447 -56 451
rect -93 443 -79 447
rect -65 443 -56 447
rect -121 435 -113 439
rect -139 328 -135 423
rect -121 415 -117 435
rect -93 427 -85 431
rect -82 431 -79 443
rect -82 427 -75 431
rect -88 423 -85 427
rect -88 419 -75 423
rect -60 415 -56 443
rect -53 443 -49 463
rect -121 411 -113 415
rect -65 411 -60 415
rect -121 380 -117 411
rect -82 388 -78 393
rect -93 384 -75 388
rect -121 376 -113 380
rect -37 380 -33 475
rect -29 569 -25 590
rect -29 454 -25 564
rect -21 497 -17 547
rect -21 442 -17 492
rect -13 513 -9 664
rect 12 651 16 664
rect 44 651 48 665
rect 63 664 67 668
rect 71 664 156 668
rect 12 647 20 651
rect 44 647 52 651
rect 4 643 5 647
rect 12 641 16 647
rect 44 641 48 647
rect 39 637 48 641
rect 4 631 5 635
rect 12 631 16 637
rect 152 631 156 664
rect 12 627 20 631
rect 62 627 66 631
rect 70 627 156 631
rect 2 601 81 605
rect 2 577 6 601
rect 77 598 81 601
rect 72 594 95 598
rect 10 589 49 593
rect 1 561 5 564
rect 10 552 14 589
rect 74 585 77 589
rect 103 585 119 589
rect 26 577 34 581
rect 6 548 14 552
rect 18 540 22 565
rect 26 565 30 577
rect 86 573 90 577
rect 74 569 90 573
rect 26 561 34 565
rect 26 548 30 561
rect 74 552 77 556
rect 86 548 90 569
rect 115 565 119 585
rect 152 565 156 627
rect 111 561 115 565
rect 119 561 128 565
rect 132 561 156 565
rect 26 544 34 548
rect 86 544 91 548
rect 18 536 89 540
rect 85 532 89 536
rect 74 528 93 532
rect 14 524 49 528
rect 74 519 77 523
rect 115 523 119 561
rect 103 519 119 523
rect 70 513 74 519
rect -13 509 70 513
rect -13 474 -9 509
rect 44 482 48 485
rect 39 478 55 482
rect -13 470 13 474
rect 17 470 21 474
rect 152 474 156 561
rect -121 372 -117 376
rect -84 372 -80 377
rect -65 376 -33 380
rect -121 368 -113 372
rect -89 369 -75 372
rect -121 356 -117 368
rect -89 364 -86 369
rect -93 360 -86 364
rect -121 352 -113 356
rect -60 356 -56 376
rect -128 328 -124 340
rect -139 324 -128 328
rect -121 340 -117 352
rect -83 348 -79 353
rect -65 352 -56 356
rect -60 348 -56 352
rect -93 344 -79 348
rect -65 344 -56 348
rect -121 336 -113 340
rect -139 230 -135 324
rect -121 316 -117 336
rect -93 328 -85 332
rect -82 332 -79 344
rect -82 328 -75 332
rect -88 324 -85 328
rect -88 320 -75 324
rect -60 316 -56 344
rect -53 344 -49 364
rect -121 312 -113 316
rect -65 312 -60 316
rect -121 282 -117 312
rect -82 290 -78 295
rect -93 286 -75 290
rect -121 278 -113 282
rect -37 282 -33 376
rect -121 274 -117 278
rect -84 274 -80 279
rect -65 278 -33 282
rect -121 270 -113 274
rect -89 271 -75 274
rect -121 258 -117 270
rect -89 266 -86 271
rect -93 262 -86 266
rect -121 254 -113 258
rect -60 258 -56 278
rect -128 230 -124 242
rect -139 226 -128 230
rect -121 242 -117 254
rect -83 250 -79 255
rect -65 254 -56 258
rect -60 250 -56 254
rect -93 246 -79 250
rect -65 246 -56 250
rect -121 238 -113 242
rect -139 133 -135 226
rect -121 218 -117 238
rect -93 230 -85 234
rect -82 234 -79 246
rect -82 230 -75 234
rect -88 226 -85 230
rect -88 222 -75 226
rect -60 218 -56 246
rect -53 246 -49 266
rect -121 214 -113 218
rect -65 214 -60 218
rect -121 185 -117 214
rect -82 193 -78 198
rect -93 189 -75 193
rect -121 181 -113 185
rect -37 185 -33 278
rect -29 371 -25 393
rect -29 257 -25 366
rect -21 300 -17 350
rect -21 245 -17 295
rect -13 315 -9 470
rect 12 457 16 470
rect 44 457 48 471
rect 63 470 67 474
rect 71 470 156 474
rect 12 453 20 457
rect 44 453 52 457
rect 4 449 5 453
rect 12 447 16 453
rect 44 447 48 453
rect 39 443 48 447
rect 4 437 5 441
rect 12 437 16 443
rect 152 437 156 470
rect 12 433 20 437
rect 62 433 66 437
rect 70 433 156 437
rect 2 403 81 407
rect 2 379 6 403
rect 77 400 81 403
rect 72 396 95 400
rect 10 391 49 395
rect 1 363 5 366
rect 10 354 14 391
rect 74 387 77 391
rect 103 387 119 391
rect 26 379 34 383
rect 6 350 14 354
rect 18 342 22 367
rect 26 367 30 379
rect 86 375 90 379
rect 74 371 90 375
rect 26 363 34 367
rect 26 350 30 363
rect 74 354 77 358
rect 86 350 90 371
rect 115 367 119 387
rect 152 367 156 433
rect 111 363 115 367
rect 119 363 128 367
rect 132 363 156 367
rect 26 346 34 350
rect 86 346 91 350
rect 18 338 89 342
rect 85 334 89 338
rect 74 330 93 334
rect 14 326 49 330
rect 74 321 77 325
rect 115 325 119 363
rect 103 321 119 325
rect 70 315 74 321
rect -13 311 70 315
rect -13 277 -9 311
rect 44 285 48 288
rect 39 281 55 285
rect -13 273 13 277
rect 17 273 21 277
rect 152 277 156 363
rect -121 177 -117 181
rect -84 177 -80 182
rect -65 181 -33 185
rect -121 173 -113 177
rect -89 174 -75 177
rect -121 161 -117 173
rect -89 169 -86 174
rect -93 165 -86 169
rect -121 157 -113 161
rect -60 161 -56 181
rect -128 133 -124 145
rect -139 129 -128 133
rect -121 145 -117 157
rect -83 153 -79 158
rect -65 157 -56 161
rect -60 153 -56 157
rect -93 149 -79 153
rect -65 149 -56 153
rect -121 141 -113 145
rect -139 34 -135 129
rect -121 121 -117 141
rect -93 133 -85 137
rect -82 137 -79 149
rect -82 133 -75 137
rect -88 129 -85 133
rect -88 125 -75 129
rect -60 121 -56 149
rect -53 149 -49 169
rect -121 117 -113 121
rect -65 117 -60 121
rect -121 85 -117 117
rect -82 93 -78 98
rect -93 89 -75 93
rect -121 81 -113 85
rect -37 85 -33 181
rect -121 77 -117 81
rect -84 77 -80 82
rect -65 81 -33 85
rect -121 73 -113 77
rect -89 74 -75 77
rect -121 61 -117 73
rect -89 69 -86 74
rect -93 65 -86 69
rect -121 57 -113 61
rect -60 61 -56 81
rect -128 33 -124 45
rect -134 29 -128 33
rect -121 45 -117 57
rect -83 53 -79 58
rect -65 57 -56 61
rect -60 53 -56 57
rect -93 49 -79 53
rect -65 49 -56 53
rect -121 41 -113 45
rect -121 21 -117 41
rect -93 33 -85 37
rect -82 37 -79 49
rect -82 33 -75 37
rect -88 29 -85 33
rect -88 25 -75 29
rect -60 21 -56 49
rect -53 49 -49 69
rect -121 17 -113 21
rect -65 17 -60 21
rect -37 -5 -33 81
rect -29 168 -25 198
rect -29 42 -25 163
rect -21 103 -17 147
rect -21 30 -17 98
rect -13 112 -9 273
rect 12 260 16 273
rect 44 260 48 274
rect 63 273 67 277
rect 71 273 156 277
rect 12 256 20 260
rect 44 256 52 260
rect 4 252 5 256
rect 12 250 16 256
rect 44 250 48 256
rect 39 246 48 250
rect 4 240 5 244
rect 12 240 16 246
rect 152 240 156 273
rect 12 236 20 240
rect 62 236 66 240
rect 70 236 156 240
rect 2 200 81 204
rect 2 176 6 200
rect 77 197 81 200
rect 72 193 95 197
rect 10 188 49 192
rect 1 160 5 163
rect 10 151 14 188
rect 74 184 77 188
rect 103 184 119 188
rect 26 176 34 180
rect 6 147 14 151
rect 18 139 22 164
rect 26 164 30 176
rect 86 172 90 176
rect 74 168 90 172
rect 26 160 34 164
rect 26 147 30 160
rect 74 151 77 155
rect 86 147 90 168
rect 115 164 119 184
rect 152 164 156 236
rect 111 160 115 164
rect 119 160 128 164
rect 132 160 156 164
rect 26 143 34 147
rect 86 143 91 147
rect 18 135 89 139
rect 85 131 89 135
rect 74 127 93 131
rect 14 123 49 127
rect 74 118 77 122
rect 115 122 119 160
rect 103 118 119 122
rect 70 112 74 118
rect -13 108 70 112
rect -13 62 -9 108
rect 44 70 48 73
rect 39 66 55 70
rect -13 58 13 62
rect 17 58 21 62
rect 152 62 156 160
rect 160 851 164 1025
rect 168 887 172 1025
rect 160 723 164 846
rect 168 733 172 882
rect 176 861 180 1025
rect 184 897 188 1025
rect 160 504 164 718
rect 168 513 172 728
rect 176 713 180 856
rect 160 284 164 499
rect 168 304 172 508
rect 176 489 180 708
rect 184 687 188 892
rect 192 871 196 1025
rect 200 933 204 1025
rect 192 697 196 866
rect 176 407 180 484
rect 184 469 188 682
rect 192 609 196 692
rect 200 661 204 928
rect 208 907 212 1025
rect 216 943 220 1025
rect 224 1002 228 1025
rect 224 917 228 997
rect 232 964 236 1030
rect 320 972 324 975
rect 315 968 331 972
rect 374 969 378 1030
rect 461 994 465 1004
rect 450 990 468 994
rect 422 982 430 986
rect 422 978 426 982
rect 459 978 463 983
rect 478 982 538 986
rect 422 974 430 978
rect 454 975 468 978
rect 422 969 426 974
rect 454 970 457 975
rect 374 965 426 969
rect 450 966 457 970
rect 232 960 289 964
rect 293 960 297 964
rect 208 807 212 902
rect 224 829 228 912
rect 232 842 236 960
rect 320 946 324 961
rect 339 960 343 964
rect 347 960 370 964
rect 314 942 328 946
rect 257 938 259 942
rect 257 928 259 932
rect 274 920 278 933
rect 257 912 259 916
rect 266 907 274 911
rect 257 902 259 906
rect 257 892 259 896
rect 257 882 259 886
rect 257 866 259 870
rect 266 865 270 907
rect 310 901 314 924
rect 322 920 326 942
rect 348 933 356 937
rect 322 916 328 920
rect 344 911 348 924
rect 274 874 278 887
rect 266 861 274 865
rect 257 856 259 860
rect 257 846 259 850
rect 266 846 270 861
rect 310 855 314 878
rect 328 874 332 897
rect 352 891 356 933
rect 348 887 356 891
rect 344 865 348 878
rect 352 846 356 887
rect 366 846 370 960
rect 270 842 274 846
rect 348 842 352 846
rect 356 842 370 846
rect 232 838 270 842
rect 208 671 212 802
rect 232 754 236 838
rect 320 762 324 765
rect 315 758 331 762
rect 232 750 289 754
rect 293 750 297 754
rect 366 754 370 842
rect 208 635 212 666
rect 232 652 236 750
rect 266 732 274 736
rect 257 728 259 732
rect 257 718 259 722
rect 257 708 259 712
rect 257 692 259 696
rect 266 691 270 732
rect 274 708 278 723
rect 320 717 324 751
rect 339 750 343 754
rect 347 750 370 754
rect 314 713 324 717
rect 320 700 324 713
rect 314 696 324 700
rect 328 708 332 732
rect 348 723 356 727
rect 328 700 332 704
rect 266 687 274 691
rect 257 682 259 686
rect 257 666 259 670
rect 274 665 278 678
rect 320 674 324 696
rect 314 670 324 674
rect 328 674 332 687
rect 352 682 356 723
rect 348 678 356 682
rect 320 665 324 670
rect 320 661 328 665
rect 352 664 356 678
rect 257 656 259 660
rect 352 656 356 660
rect 366 656 370 750
rect 270 652 274 656
rect 348 652 370 656
rect 232 648 270 652
rect 192 479 196 604
rect 232 533 236 648
rect 321 541 325 544
rect 316 537 332 541
rect 232 529 290 533
rect 294 529 298 533
rect 366 533 370 652
rect 192 422 196 474
rect 232 460 236 529
rect 257 508 260 512
rect 257 500 260 504
rect 276 492 280 504
rect 321 500 325 530
rect 340 529 344 533
rect 348 529 370 533
rect 316 496 325 500
rect 257 484 260 488
rect 321 483 325 496
rect 316 479 325 483
rect 330 483 334 512
rect 350 504 358 508
rect 346 492 350 496
rect 257 474 260 478
rect 321 473 325 479
rect 321 469 330 473
rect 354 468 358 504
rect 257 464 260 468
rect 366 464 370 529
rect 272 460 276 464
rect 350 460 370 464
rect 232 456 272 460
rect 176 294 180 402
rect 232 328 236 456
rect 321 336 325 339
rect 316 332 332 336
rect 232 324 290 328
rect 294 324 298 328
rect 366 328 370 460
rect 160 252 164 279
rect 176 268 180 289
rect 232 275 236 324
rect 321 307 325 325
rect 340 324 344 328
rect 348 324 370 328
rect 366 307 370 324
rect 319 303 332 307
rect 353 303 370 307
rect 257 299 264 303
rect 328 298 332 303
rect 319 294 324 298
rect 328 294 333 298
rect 257 289 264 293
rect 275 284 279 288
rect 257 279 264 283
rect 271 275 275 284
rect 320 279 324 294
rect 357 288 361 303
rect 357 279 361 284
rect 319 275 324 279
rect 353 275 361 279
rect 232 271 275 275
rect 160 78 164 247
rect 12 45 16 58
rect 44 45 48 59
rect 63 58 67 62
rect 71 58 156 62
rect 12 41 20 45
rect 44 41 52 45
rect 4 37 5 41
rect 12 35 16 41
rect 44 35 48 41
rect 39 31 48 35
rect 4 25 5 29
rect 12 25 16 31
rect 152 25 156 58
rect 12 21 20 25
rect 62 21 66 25
rect 70 21 156 25
rect 152 -5 156 21
rect 366 -5 370 303
rect 374 773 378 965
rect 422 962 426 965
rect 422 958 430 962
rect 483 962 487 982
rect 415 934 419 946
rect 398 930 415 934
rect 422 946 426 958
rect 460 954 464 959
rect 478 958 487 962
rect 483 954 487 958
rect 450 950 464 954
rect 478 950 487 954
rect 422 942 430 946
rect 398 884 402 930
rect 422 922 426 942
rect 450 934 458 938
rect 461 938 464 950
rect 461 934 468 938
rect 455 930 458 934
rect 455 926 468 930
rect 483 922 487 950
rect 490 950 494 970
rect 422 918 430 922
rect 478 918 483 922
rect 397 861 476 865
rect 397 837 401 861
rect 472 858 476 861
rect 467 854 490 858
rect 405 849 444 853
rect 396 821 400 824
rect 405 812 409 849
rect 469 845 472 849
rect 498 845 514 849
rect 421 837 429 841
rect 396 808 397 812
rect 401 808 409 812
rect 413 800 417 825
rect 421 825 425 837
rect 481 833 485 837
rect 469 829 485 833
rect 421 821 429 825
rect 421 808 425 821
rect 469 812 472 816
rect 481 808 485 829
rect 510 825 514 845
rect 534 825 538 982
rect 577 931 581 1030
rect 616 939 620 949
rect 605 935 623 939
rect 577 927 585 931
rect 577 923 581 927
rect 614 923 618 928
rect 633 927 658 931
rect 577 919 585 923
rect 609 920 623 923
rect 577 907 581 919
rect 609 915 612 920
rect 605 911 612 915
rect 577 903 585 907
rect 638 907 642 927
rect 506 821 510 825
rect 514 821 523 825
rect 527 821 538 825
rect 421 804 429 808
rect 481 804 486 808
rect 413 796 484 800
rect 480 792 484 796
rect 469 788 488 792
rect 409 784 444 788
rect 469 779 472 783
rect 510 783 514 821
rect 498 779 514 783
rect 465 773 469 779
rect 374 769 465 773
rect 374 579 378 769
rect 397 667 476 671
rect 397 643 401 667
rect 472 664 476 667
rect 467 660 490 664
rect 405 655 444 659
rect 396 627 400 630
rect 405 618 409 655
rect 469 651 472 655
rect 498 651 514 655
rect 421 643 429 647
rect 396 614 397 618
rect 401 614 409 618
rect 413 606 417 631
rect 421 631 425 643
rect 481 639 485 643
rect 469 635 485 639
rect 421 627 429 631
rect 421 614 425 627
rect 469 618 472 622
rect 481 614 485 635
rect 510 631 514 651
rect 534 631 538 821
rect 506 627 510 631
rect 514 627 523 631
rect 527 627 538 631
rect 421 610 429 614
rect 481 610 486 614
rect 413 602 484 606
rect 480 598 484 602
rect 469 594 488 598
rect 409 590 444 594
rect 469 585 472 589
rect 510 589 514 627
rect 498 585 514 589
rect 465 579 469 585
rect 374 575 465 579
rect 374 366 378 575
rect 397 454 476 458
rect 397 430 401 454
rect 472 451 476 454
rect 467 447 490 451
rect 405 442 444 446
rect 396 414 400 417
rect 405 405 409 442
rect 469 438 472 442
rect 498 438 514 442
rect 421 430 429 434
rect 396 401 397 405
rect 401 401 409 405
rect 413 393 417 418
rect 421 418 425 430
rect 481 426 485 430
rect 469 422 485 426
rect 421 414 429 418
rect 421 401 425 414
rect 469 405 472 409
rect 481 401 485 422
rect 510 418 514 438
rect 534 418 538 627
rect 506 414 510 418
rect 514 414 523 418
rect 527 414 538 418
rect 421 397 429 401
rect 481 397 486 401
rect 413 389 484 393
rect 480 385 484 389
rect 469 381 488 385
rect 409 377 444 381
rect 469 372 472 376
rect 510 376 514 414
rect 498 372 514 376
rect 465 366 469 372
rect 374 362 465 366
rect 374 212 378 362
rect 397 300 476 304
rect 397 276 401 300
rect 472 297 476 300
rect 467 293 490 297
rect 405 288 444 292
rect 396 260 400 263
rect 405 251 409 288
rect 469 284 472 288
rect 498 284 514 288
rect 421 276 429 280
rect 396 247 397 251
rect 401 247 409 251
rect 413 239 417 264
rect 421 264 425 276
rect 481 272 485 276
rect 469 268 485 272
rect 421 260 429 264
rect 421 247 425 260
rect 469 251 472 255
rect 481 247 485 268
rect 510 264 514 284
rect 534 264 538 414
rect 506 260 510 264
rect 514 260 523 264
rect 527 260 538 264
rect 421 243 429 247
rect 481 243 486 247
rect 413 235 484 239
rect 480 231 484 235
rect 469 227 488 231
rect 409 223 444 227
rect 469 218 472 222
rect 510 222 514 260
rect 498 218 514 222
rect 465 212 469 218
rect 374 208 465 212
rect 534 -5 538 260
rect 570 879 574 891
rect 542 875 570 879
rect 577 891 581 903
rect 615 899 619 904
rect 633 903 642 907
rect 638 899 642 903
rect 605 895 619 899
rect 633 895 642 899
rect 577 887 585 891
rect 542 685 546 875
rect 577 867 581 887
rect 605 879 613 883
rect 616 883 619 895
rect 616 879 623 883
rect 610 875 613 879
rect 610 871 623 875
rect 638 867 642 895
rect 645 895 649 915
rect 577 863 585 867
rect 633 863 638 867
rect 577 737 581 863
rect 616 745 620 755
rect 605 741 623 745
rect 577 733 585 737
rect 654 737 658 927
rect 577 729 581 733
rect 614 729 618 734
rect 633 733 658 737
rect 577 725 585 729
rect 609 726 623 729
rect 577 713 581 725
rect 609 721 612 726
rect 605 717 612 721
rect 577 709 585 713
rect 638 713 642 733
rect 570 685 574 697
rect 542 681 570 685
rect 577 697 581 709
rect 615 705 619 710
rect 633 709 642 713
rect 638 705 642 709
rect 605 701 619 705
rect 633 701 642 705
rect 577 693 585 697
rect 542 472 546 681
rect 577 673 581 693
rect 605 685 613 689
rect 616 689 619 701
rect 616 685 623 689
rect 610 681 613 685
rect 610 677 623 681
rect 638 673 642 701
rect 645 701 649 721
rect 577 669 585 673
rect 633 669 638 673
rect 577 524 581 669
rect 616 532 620 542
rect 605 528 623 532
rect 577 520 585 524
rect 654 524 658 733
rect 577 516 581 520
rect 614 516 618 521
rect 633 520 658 524
rect 577 512 585 516
rect 609 513 623 516
rect 577 500 581 512
rect 609 508 612 513
rect 605 504 612 508
rect 577 496 585 500
rect 638 500 642 520
rect 570 472 574 484
rect 542 468 570 472
rect 577 484 581 496
rect 615 492 619 497
rect 633 496 642 500
rect 638 492 642 496
rect 605 488 619 492
rect 633 488 642 492
rect 577 480 585 484
rect 542 318 546 468
rect 577 460 581 480
rect 605 472 613 476
rect 616 476 619 488
rect 616 472 623 476
rect 610 468 613 472
rect 610 464 623 468
rect 638 460 642 488
rect 645 488 649 508
rect 577 456 585 460
rect 633 456 638 460
rect 577 370 581 456
rect 616 378 620 388
rect 605 374 623 378
rect 577 366 585 370
rect 654 370 658 520
rect 577 362 581 366
rect 614 362 618 367
rect 633 366 658 370
rect 577 358 585 362
rect 609 359 623 362
rect 577 346 581 358
rect 609 354 612 359
rect 605 350 612 354
rect 577 342 585 346
rect 638 346 642 366
rect 570 318 574 330
rect 542 314 570 318
rect 577 330 581 342
rect 615 338 619 343
rect 633 342 642 346
rect 638 338 642 342
rect 605 334 619 338
rect 633 334 642 338
rect 577 326 585 330
rect 542 210 546 314
rect 577 306 581 326
rect 605 318 613 322
rect 616 322 619 334
rect 616 318 623 322
rect 610 314 613 318
rect 610 310 623 314
rect 638 306 642 334
rect 645 334 649 354
rect 577 302 585 306
rect 633 302 638 306
rect 577 262 581 302
rect 616 270 620 280
rect 605 266 623 270
rect 577 258 585 262
rect 654 262 658 366
rect 577 254 581 258
rect 614 254 618 259
rect 633 258 658 262
rect 577 250 585 254
rect 609 251 623 254
rect 577 238 581 250
rect 609 246 612 251
rect 605 242 612 246
rect 577 234 585 238
rect 638 238 642 258
rect 570 210 574 222
rect 542 206 570 210
rect 577 222 581 234
rect 615 230 619 235
rect 633 234 642 238
rect 638 230 642 234
rect 605 226 619 230
rect 633 226 642 230
rect 577 218 585 222
rect 542 9 546 206
rect 577 198 581 218
rect 605 210 613 214
rect 616 214 619 226
rect 616 210 623 214
rect 610 206 613 210
rect 610 202 623 206
rect 638 198 642 226
rect 645 226 649 246
rect 577 194 585 198
rect 633 194 638 198
rect 654 -5 658 258
rect -37 -9 658 -5
<< m2contact >>
rect -82 986 -77 991
rect -29 986 -24 991
rect -82 886 -77 891
rect -82 786 -77 791
rect -29 957 -24 962
rect -21 941 -16 946
rect -22 886 -17 891
rect -29 843 -24 848
rect 0 957 5 962
rect -3 941 2 946
rect 77 977 82 982
rect 86 970 91 975
rect 77 945 82 950
rect 9 917 14 922
rect 77 912 82 917
rect 44 879 49 884
rect -21 831 -16 836
rect -82 686 -77 691
rect -82 590 -77 595
rect -29 786 -24 791
rect -29 762 -24 767
rect -21 746 -16 751
rect -22 686 -17 691
rect -29 643 -24 648
rect -1 843 4 848
rect -1 831 4 836
rect 0 762 5 767
rect -3 746 2 751
rect 77 782 82 787
rect 86 775 91 780
rect 77 750 82 755
rect 9 722 14 727
rect 77 717 82 722
rect 44 679 49 684
rect -21 631 -16 636
rect -82 492 -77 497
rect -82 393 -77 398
rect -29 590 -24 595
rect -29 564 -24 569
rect -21 547 -16 552
rect -22 492 -17 497
rect -29 449 -24 454
rect -1 643 4 648
rect -1 631 4 636
rect 0 564 5 569
rect 77 584 82 589
rect 86 577 91 582
rect -3 547 2 552
rect 77 552 82 557
rect 9 524 14 529
rect 77 519 82 524
rect 44 485 49 490
rect -21 437 -16 442
rect -82 295 -77 300
rect -82 198 -77 203
rect -29 393 -24 398
rect -29 366 -24 371
rect -21 350 -16 355
rect -22 295 -17 300
rect -29 252 -24 257
rect -1 449 4 454
rect -1 437 4 442
rect 0 366 5 371
rect -3 350 2 355
rect 77 386 82 391
rect 86 379 91 384
rect 77 354 82 359
rect 9 326 14 331
rect 77 321 82 326
rect 44 288 49 293
rect -21 240 -16 245
rect -82 98 -77 103
rect -139 29 -134 34
rect -29 198 -24 203
rect -29 163 -24 168
rect -21 147 -16 152
rect -22 98 -17 103
rect -29 37 -24 42
rect -1 252 4 257
rect -1 240 4 245
rect 0 163 5 168
rect -3 147 2 152
rect 77 183 82 188
rect 86 176 91 181
rect 77 151 82 156
rect 9 123 14 128
rect 77 118 82 123
rect 44 73 49 78
rect 168 882 173 887
rect 160 846 165 851
rect 184 892 189 897
rect 176 856 181 861
rect 168 728 173 733
rect 160 718 165 723
rect 176 708 181 713
rect 168 508 173 513
rect 160 499 165 504
rect 200 928 205 933
rect 192 866 197 871
rect 192 692 197 697
rect 184 682 189 687
rect 176 484 181 489
rect 223 997 228 1002
rect 216 938 221 943
rect 320 975 325 980
rect 224 912 229 917
rect 208 902 213 907
rect 252 938 257 943
rect 252 928 257 933
rect 252 912 257 917
rect 252 902 257 907
rect 252 892 257 897
rect 252 882 257 887
rect 252 866 257 871
rect 252 856 257 861
rect 252 846 257 851
rect 224 824 229 829
rect 207 802 212 807
rect 320 765 325 770
rect 208 666 213 671
rect 200 656 205 661
rect 252 728 257 733
rect 252 718 257 723
rect 252 708 257 713
rect 252 692 257 697
rect 252 682 257 687
rect 252 666 257 671
rect 252 656 257 661
rect 208 630 213 635
rect 191 604 196 609
rect 321 544 326 549
rect 192 474 197 479
rect 184 464 189 469
rect 252 508 257 513
rect 252 499 257 504
rect 252 484 257 489
rect 252 474 257 479
rect 252 464 257 469
rect 192 417 197 422
rect 175 402 180 407
rect 168 299 173 304
rect 321 339 326 344
rect 176 289 181 294
rect 160 279 165 284
rect 252 299 257 304
rect 252 289 257 294
rect 252 279 257 284
rect 176 263 181 268
rect 160 247 165 252
rect 159 73 164 78
rect -1 37 4 42
rect -21 25 -16 30
rect -1 25 4 30
rect 410 922 415 927
rect 398 879 403 884
rect 395 824 400 829
rect 391 808 396 813
rect 472 844 477 849
rect 481 837 486 842
rect 472 812 477 817
rect 404 784 409 789
rect 472 779 477 784
rect 395 630 400 635
rect 391 614 396 619
rect 472 650 477 655
rect 481 643 486 648
rect 472 618 477 623
rect 404 590 409 595
rect 472 585 477 590
rect 395 417 400 422
rect 391 401 396 406
rect 472 437 477 442
rect 481 430 486 435
rect 472 405 477 410
rect 404 377 409 382
rect 472 372 477 377
rect 395 263 400 268
rect 391 247 396 252
rect 472 283 477 288
rect 481 276 486 281
rect 472 251 477 256
rect 404 223 409 228
rect 472 218 477 223
rect 542 879 547 884
rect 565 867 570 872
rect 565 673 570 678
rect 565 460 570 465
rect 565 306 570 311
rect 565 198 570 203
rect 542 4 547 9
<< pdm12contact >>
rect 276 512 281 517
rect 276 469 281 474
<< metal2 >>
rect 86 997 223 1002
rect -77 986 -29 991
rect -24 957 0 962
rect 5 958 14 962
rect -16 941 -3 946
rect 9 922 14 958
rect 78 950 82 977
rect 86 975 91 997
rect 325 975 409 980
rect 78 917 82 945
rect 141 938 216 943
rect 221 938 252 943
rect -77 886 -22 891
rect 141 884 146 938
rect 205 928 252 933
rect 404 927 409 975
rect 404 922 410 927
rect 229 912 252 917
rect 213 902 252 907
rect 189 892 252 897
rect 49 879 146 884
rect 173 882 252 887
rect 403 879 542 884
rect 197 866 252 871
rect 481 867 565 872
rect 181 856 252 861
rect -24 843 -1 848
rect 165 846 252 851
rect -16 831 -1 836
rect 229 824 395 829
rect 400 825 409 829
rect 320 808 391 813
rect 86 802 207 807
rect -77 786 -29 791
rect -24 762 0 767
rect 5 763 14 767
rect -16 746 -3 751
rect 9 727 14 763
rect 78 755 82 782
rect 86 780 91 802
rect 320 770 325 808
rect 404 789 409 825
rect 473 817 477 844
rect 481 842 486 867
rect 473 784 477 812
rect 78 722 82 750
rect 173 728 252 733
rect 165 718 252 723
rect 181 708 252 713
rect 197 692 252 697
rect -77 686 -22 691
rect 49 679 95 684
rect 189 682 252 687
rect 90 661 95 679
rect 481 673 565 678
rect 213 666 252 671
rect 90 656 200 661
rect 205 656 252 661
rect -24 643 -1 648
rect -16 631 -1 636
rect 213 630 395 635
rect 400 631 409 635
rect 321 614 391 619
rect 86 604 191 609
rect -77 590 -29 595
rect -24 564 0 569
rect 5 565 14 569
rect -16 547 -3 552
rect 9 529 14 565
rect 78 557 82 584
rect 86 582 91 604
rect 78 524 82 552
rect 321 549 326 614
rect 404 595 409 631
rect 473 623 477 650
rect 481 648 486 673
rect 473 590 477 618
rect 173 508 252 513
rect 269 512 276 517
rect 165 499 252 504
rect -77 492 -22 497
rect 49 485 115 490
rect 110 469 115 485
rect 181 484 252 489
rect 197 474 252 479
rect 269 474 274 512
rect 269 469 276 474
rect 110 464 184 469
rect 189 464 252 469
rect 481 460 565 465
rect -24 449 -1 454
rect -16 437 -1 442
rect 197 417 395 422
rect 400 418 409 422
rect 86 402 175 407
rect -77 393 -29 398
rect -24 366 0 371
rect 5 367 14 371
rect -16 350 -3 355
rect 9 331 14 367
rect 78 359 82 386
rect 86 384 91 402
rect 321 401 391 406
rect 78 326 82 354
rect 321 344 326 401
rect 404 382 409 418
rect 473 410 477 437
rect 481 435 486 460
rect 473 377 477 405
rect 481 306 565 311
rect -77 295 -22 300
rect 44 299 168 304
rect 173 299 252 304
rect 44 293 49 299
rect 181 289 252 294
rect 165 279 252 284
rect 181 263 395 268
rect 400 264 409 268
rect -24 252 -1 257
rect 165 247 391 252
rect -16 240 -1 245
rect 404 228 409 264
rect 473 256 477 283
rect 481 281 486 306
rect 473 223 477 251
rect -77 198 -29 203
rect 86 198 565 203
rect -24 163 0 168
rect 5 163 14 168
rect -16 147 -3 152
rect 9 128 14 163
rect 78 156 82 183
rect 86 181 91 198
rect 78 123 82 151
rect -77 98 -22 103
rect 49 73 159 78
rect -24 37 -1 42
rect -139 4 -134 29
rect -16 25 -1 30
rect -139 -1 547 4
<< labels >>
rlabel metal1 161 1024 163 1025 5 G0
rlabel metal1 169 1024 171 1025 5 G1
rlabel metal1 177 1024 179 1025 5 P1
rlabel metal1 185 1024 187 1025 5 G2
rlabel metal1 193 1024 195 1025 5 P2
rlabel metal1 201 1024 203 1025 5 G3
rlabel metal1 209 1024 211 1025 5 P3
rlabel metal1 217 1024 219 1025 5 G4
rlabel metal1 225 1024 227 1025 5 P4
rlabel metal1 321 953 323 954 7 C5_bar
rlabel metal1 342 960 343 964 7 gnd
rlabel metal1 294 960 295 964 7 vdd
rlabel polycontact 259 939 260 941 7 G4
rlabel polycontact 259 929 260 931 7 G3
rlabel polycontact 259 913 260 915 7 P4
rlabel polycontact 259 903 260 905 7 P3
rlabel polycontact 259 893 260 895 7 G2
rlabel polycontact 259 883 260 885 7 G1
rlabel polycontact 259 867 260 869 7 P2
rlabel polycontact 259 857 260 859 7 P1
rlabel polycontact 259 847 260 849 7 G0
rlabel psubstratepcontact 352 842 356 846 7 gnd
rlabel nsubstratencontact 267 843 268 845 7 vdd
rlabel metal1 321 743 323 744 7 C4_bar
rlabel metal1 342 750 343 754 7 gnd
rlabel metal1 294 750 295 754 7 vdd
rlabel polycontact 259 729 260 731 3 G1
rlabel polycontact 259 719 260 721 3 G0
rlabel polycontact 259 709 260 711 3 P1
rlabel polycontact 259 693 260 695 3 P2
rlabel polycontact 259 683 260 685 3 G2
rlabel polycontact 259 667 260 669 3 P3
rlabel polycontact 259 657 260 659 3 G3
rlabel nsubstratencontact 267 653 269 655 7 vdd
rlabel metal1 353 652 355 655 8 gnd
rlabel metal1 322 522 324 523 7 C3_bar
rlabel metal1 343 529 344 533 7 gnd
rlabel metal1 295 529 296 533 7 vdd
rlabel metal1 258 509 259 511 3 G1
rlabel metal1 258 501 259 503 3 G0
rlabel metal1 258 485 259 487 3 P1
rlabel metal1 258 475 259 477 3 P2
rlabel metal1 258 465 259 467 3 G2
rlabel nsubstratencontact 271 461 272 463 7 vdd
rlabel metal1 355 460 356 462 7 gnd
rlabel metal1 271 284 272 287 3 vdd
rlabel metal1 262 279 263 282 3 G0
rlabel metal1 262 299 263 302 3 G1
rlabel metal1 295 324 296 328 7 vdd
rlabel metal1 343 324 344 328 7 gnd
rlabel metal1 323 311 324 316 7 C2_bar
rlabel metal1 358 275 359 278 8 gnd
rlabel metal1 262 289 263 292 3 P1
rlabel polycontact 1 950 5 954 1 B4
rlabel polycontact 2 941 6 945 1 A4
rlabel metal1 106 978 107 982 7 gnd
rlabel nsubstratencontact 70 902 74 906 1 vdd
rlabel metal1 46 854 47 859 1 G4_bar
rlabel m2contact 1 844 2 846 1 B4
rlabel m2contact 1 832 2 834 1 A4
rlabel metal1 66 864 67 868 7 gnd
rlabel metal1 18 864 19 868 7 vdd
rlabel metal1 12 827 13 831 3 vdd
rlabel metal1 64 827 66 828 8 gnd
rlabel polycontact 1 755 5 759 1 B3
rlabel polycontact 2 746 6 750 1 A3
rlabel metal1 113 759 119 763 7 gnd
rlabel metal1 106 783 107 787 7 gnd
rlabel nsubstratencontact 70 707 74 711 1 vdd
rlabel metal1 46 654 47 659 1 G3_bar
rlabel m2contact 1 632 2 634 1 A3
rlabel metal1 66 664 67 668 7 gnd
rlabel metal1 18 664 19 668 7 vdd
rlabel metal1 12 627 13 631 3 vdd
rlabel metal1 64 627 66 628 8 gnd
rlabel nsubstratencontact 70 509 74 513 1 vdd
rlabel metal1 106 585 107 589 7 gnd
rlabel metal1 113 561 119 565 7 gnd
rlabel polycontact 2 548 6 552 3 A2
rlabel polycontact 1 557 5 561 3 B2
rlabel metal1 64 433 66 434 8 gnd
rlabel metal1 12 433 13 437 3 vdd
rlabel metal1 18 470 19 474 7 vdd
rlabel metal1 66 470 67 474 7 gnd
rlabel m2contact 1 438 2 440 1 A2
rlabel m2contact 1 450 2 452 1 B2
rlabel metal1 46 460 47 465 1 G2_bar
rlabel polycontact 1 359 5 363 3 B1
rlabel polycontact 2 350 6 354 3 A1
rlabel nsubstratencontact 70 311 74 315 1 vdd
rlabel metal1 106 387 107 391 7 gnd
rlabel metal1 113 363 119 367 7 gnd
rlabel metal1 46 263 47 268 1 G1_bar
rlabel metal1 66 273 67 277 7 gnd
rlabel metal1 18 273 19 277 7 vdd
rlabel metal1 12 236 13 240 3 vdd
rlabel metal1 64 236 66 237 8 gnd
rlabel polycontact 1 156 5 160 3 B0
rlabel nsubstratencontact 70 108 74 112 1 vdd
rlabel metal1 106 184 107 188 7 gnd
rlabel metal1 113 160 119 164 7 gnd
rlabel metal1 66 58 67 62 7 gnd
rlabel metal1 18 58 19 62 7 vdd
rlabel metal1 12 21 13 25 3 vdd
rlabel metal1 64 21 66 22 8 gnd
rlabel m2contact 1 26 2 28 1 A0
rlabel m2contact 1 38 2 40 1 B0
rlabel metal1 46 48 47 53 1 G0_bar
rlabel metal2 378 200 381 202 1 S0
rlabel polycontact 396 256 400 260 1 P1
rlabel metal1 508 260 514 264 7 gnd
rlabel metal1 501 284 502 288 7 gnd
rlabel nsubstratencontact 465 208 469 212 1 vdd
rlabel nsubstratencontact 465 362 469 366 1 vdd
rlabel metal1 501 438 502 442 7 gnd
rlabel metal1 508 414 514 418 7 gnd
rlabel metal1 508 627 514 631 7 gnd
rlabel metal1 501 651 502 655 7 gnd
rlabel nsubstratencontact 465 575 469 579 1 vdd
rlabel nsubstratencontact 465 769 469 773 1 vdd
rlabel metal1 501 845 502 849 7 gnd
rlabel metal1 508 821 514 825 7 gnd
rlabel polycontact 397 247 401 251 1 G0
rlabel polycontact 397 401 401 405 1 C2
rlabel polycontact 396 410 400 414 1 P2
rlabel polycontact 397 614 401 618 1 C3
rlabel polycontact 396 623 400 627 1 P3
rlabel polycontact 397 808 401 812 1 C4
rlabel polycontact 396 817 400 821 1 P4
rlabel metal2 484 869 487 871 1 S4
rlabel metal2 484 674 487 676 1 S3
rlabel metal2 483 461 486 463 1 S2
rlabel metal2 484 308 487 310 1 S1
rlabel polycontact -128 29 -124 33 3 CLK
rlabel polycontact -128 21 -124 25 3 A0_reg
rlabel m2contact -82 98 -78 102 1 A0
rlabel metal1 -121 68 -117 72 1 vdd
rlabel metal1 -60 51 -56 55 1 gnd
rlabel polycontact -128 121 -124 125 3 B0_reg
rlabel polycontact -128 129 -124 133 3 CLK
rlabel metal1 -82 195 -78 199 1 B0
rlabel metal1 -121 169 -117 173 1 vdd
rlabel metal1 -60 173 -56 177 1 gnd
rlabel polycontact 2 147 6 151 3 A0
rlabel polycontact -128 218 -124 222 3 A1_reg
rlabel polycontact -128 226 -124 230 3 CLK
rlabel metal1 -121 259 -117 263 1 vdd
rlabel metal1 -60 255 -56 259 1 gnd
rlabel metal1 -82 293 -78 296 1 A1
rlabel polycontact -128 316 -124 320 3 B1_reg
rlabel polycontact -128 324 -124 328 3 CLK
rlabel metal1 -121 352 -117 356 1 vdd
rlabel metal1 -60 352 -56 356 1 gnd
rlabel metal1 -82 392 -78 396 1 B1
rlabel m2contact 1 241 2 243 1 A1
rlabel m2contact 1 253 2 255 1 B1
rlabel polycontact -128 415 -124 419 3 A2_reg
rlabel polycontact -128 423 -124 427 3 CLK
rlabel metal1 -121 450 -117 454 1 vdd
rlabel metal1 -60 451 -56 455 1 gnd
rlabel metal1 -82 490 -78 494 1 A2
rlabel polycontact -128 513 -124 517 3 B2_reg
rlabel polycontact -128 521 -124 525 3 CLK
rlabel metal1 -121 545 -117 549 1 vdd
rlabel metal1 -60 545 -56 549 1 gnd
rlabel metal1 -82 588 -78 592 1 B2
rlabel m2contact 1 644 2 646 1 B3
rlabel polycontact -128 611 -124 615 3 A3_reg
rlabel polycontact -128 619 -124 623 3 CLK
rlabel metal1 -121 647 -117 651 1 vdd
rlabel metal1 -60 647 -56 651 1 gnd
rlabel metal1 -82 685 -78 689 1 A3
rlabel polycontact -128 718 -124 722 3 CLK
rlabel metal1 -82 783 -78 787 1 B3
rlabel metal1 -121 753 -117 757 1 vdd
rlabel metal1 -60 742 -56 746 1 gnd
rlabel polycontact -128 710 -124 714 3 B3_reg
rlabel polycontact -128 809 -124 813 3 A4_reg
rlabel polycontact -128 817 -124 821 3 CLK
rlabel metal1 -121 845 -117 849 1 vdd
rlabel metal1 -60 841 -56 845 1 gnd
rlabel metal1 -82 884 -78 888 1 A4
rlabel polycontact -128 906 -124 910 3 B4_reg
rlabel polycontact -128 914 -124 918 3 CLK
rlabel metal1 -121 942 -117 946 1 vdd
rlabel metal1 -60 938 -56 942 1 gnd
rlabel metal1 -82 981 -78 985 1 B4
rlabel polycontact 570 314 574 318 3 CLK
rlabel metal1 577 353 581 357 1 vdd
rlabel metal1 638 336 642 340 1 gnd
rlabel polycontact 570 206 574 210 3 CLK
rlabel metal1 577 245 581 249 1 vdd
rlabel metal1 638 228 642 232 1 gnd
rlabel polycontact 570 468 574 472 3 CLK
rlabel metal1 577 507 581 511 1 vdd
rlabel metal1 638 490 642 494 1 gnd
rlabel polycontact 570 681 574 685 3 CLK
rlabel metal1 577 720 581 724 1 vdd
rlabel metal1 638 703 642 707 1 gnd
rlabel polycontact 570 875 574 879 3 CLK
rlabel metal1 577 914 581 918 1 vdd
rlabel metal1 638 897 642 901 1 gnd
rlabel polycontact 415 930 419 934 3 CLK
rlabel metal1 422 969 426 973 1 vdd
rlabel metal1 483 952 487 956 1 gnd
rlabel polycontact 570 198 574 202 1 S0
rlabel metal1 616 275 620 279 1 Sum_out0
rlabel polycontact 570 306 574 310 1 S1
rlabel metal1 616 383 620 387 1 Sum_out1
rlabel polycontact 570 460 574 464 1 S2
rlabel metal1 616 537 620 541 1 Sum_out2
rlabel polycontact 570 673 574 677 1 S3
rlabel metal1 616 750 620 754 1 Sum_out3
rlabel polycontact 570 867 574 871 1 S4
rlabel metal1 616 943 620 947 1 Sum_out4
rlabel polycontact 415 922 419 926 1 C5
rlabel metal2 358 976 366 978 1 C5
rlabel metal1 461 998 465 1002 1 Cout_out
<< end >>
