magic
tech scmos
timestamp 1763301936
<< nwell >>
rect -21 32 26 59
rect -21 -5 57 32
rect -21 -6 23 -5
<< ntransistor >>
rect -10 -34 -8 -14
rect 0 -34 2 -14
rect 10 -34 12 -14
rect 39 -21 41 -11
<< ptransistor >>
rect -10 0 -8 40
rect 0 0 2 40
rect 10 0 12 40
rect 39 1 41 21
<< ndiffusion >>
rect -15 -30 -10 -14
rect -11 -34 -10 -30
rect -8 -34 0 -14
rect 2 -18 4 -14
rect 8 -18 10 -14
rect 2 -34 10 -18
rect 12 -30 17 -14
rect 34 -17 39 -11
rect 38 -21 39 -17
rect 41 -13 46 -11
rect 41 -17 42 -13
rect 41 -21 46 -17
rect 12 -34 13 -30
<< pdiffusion >>
rect -15 4 -10 40
rect -11 0 -10 4
rect -8 36 -6 40
rect -2 36 0 40
rect -8 0 0 36
rect 2 4 10 40
rect 2 0 4 4
rect 8 0 10 4
rect 12 4 17 40
rect 12 0 13 4
rect 38 17 39 21
rect 34 1 39 17
rect 41 7 46 21
rect 41 3 42 7
rect 41 1 46 3
<< ndcontact >>
rect -15 -34 -11 -30
rect 4 -18 8 -14
rect 34 -21 38 -17
rect 42 -17 46 -13
rect 13 -34 17 -30
<< pdcontact >>
rect -15 0 -11 4
rect -6 36 -2 40
rect 4 0 8 4
rect 13 0 17 4
rect 34 17 38 21
rect 42 3 46 7
<< psubstratepcontact >>
rect 34 -29 38 -25
rect -6 -42 -2 -38
<< nsubstratencontact >>
rect -6 44 -2 48
rect 34 25 38 29
<< polysilicon >>
rect -10 40 -8 51
rect 0 40 2 51
rect 10 40 12 51
rect 39 21 41 24
rect -10 -14 -8 0
rect 0 -14 2 0
rect 10 -14 12 0
rect 39 -11 41 1
rect 39 -24 41 -21
rect -10 -37 -8 -34
rect 0 -37 2 -34
rect 10 -37 12 -34
<< polycontact >>
rect -11 51 -7 55
rect -1 51 3 55
rect 9 51 13 55
rect 35 -6 39 -2
<< metal1 >>
rect -11 55 -7 57
rect -1 55 3 57
rect 9 55 13 57
rect -6 40 -2 44
rect 34 21 38 25
rect -15 -1 -11 0
rect 4 -1 8 0
rect -15 -5 8 -1
rect 13 -2 17 0
rect 42 -2 46 3
rect 13 -6 35 -2
rect 42 -6 53 -2
rect 13 -9 17 -6
rect 4 -13 17 -9
rect 42 -13 46 -6
rect 4 -14 8 -13
rect 34 -25 38 -21
rect -15 -38 -11 -34
rect 13 -38 17 -34
rect -15 -42 -6 -38
rect -2 -42 17 -38
<< labels >>
rlabel metal1 -6 47 -3 48 5 vdd
rlabel metal1 -11 56 -8 57 5 G0
rlabel metal1 -1 56 2 57 5 P1
rlabel metal1 9 56 12 57 5 G1
rlabel metal1 34 23 38 24 1 vdd
rlabel metal1 34 -25 38 -24 1 gnd
rlabel metal1 21 -5 26 -4 1 C2_bar
rlabel metal1 52 -5 53 -3 7 C2
rlabel metal1 -15 -40 -12 -39 2 gnd
<< end >>
