* SPICE3 file created from INV.ext - technology: scmos

.option scale=90n

M1000 Vout Vin vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1001 Vout Vin gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
C0 Vout gnd 0
C1 Vout Vin 0.0587f
C2 Vin vdd 0.03699f
C3 Vin gnd 0
C4 Vout vdd 0.01479f
C5 gnd 0 0.03709f
C6 Vout 0 0.07523f
C7 Vin 0 0.16133f
C8 vdd 0 1.18383f
