magic
tech scmos
timestamp 1763315935
<< nwell >>
rect -19 -7 79 54
rect 48 -8 79 -7
<< polysilicon >>
rect -8 40 -6 52
rect 2 40 4 52
rect 12 40 14 52
rect 28 40 30 52
rect 36 40 38 52
rect 61 18 63 21
rect -8 -14 -6 0
rect 2 -14 4 0
rect 12 -14 14 0
rect 28 -14 30 0
rect 36 -14 38 0
rect 61 -14 63 -2
rect 61 -27 63 -24
rect -8 -37 -6 -34
rect 2 -37 4 -34
rect 12 -37 14 -34
rect 28 -37 30 -34
rect 36 -37 38 -34
<< ndiffusion >>
rect -13 -30 -8 -14
rect -9 -34 -8 -30
rect -6 -18 -4 -14
rect 0 -18 2 -14
rect -6 -34 2 -18
rect 4 -18 6 -14
rect 10 -18 12 -14
rect 4 -34 12 -18
rect 14 -30 19 -14
rect 14 -34 15 -30
rect 23 -30 28 -14
rect 27 -34 28 -30
rect 30 -30 36 -14
rect 30 -34 31 -30
rect 35 -34 36 -30
rect 38 -18 39 -14
rect 38 -34 43 -18
rect 56 -20 61 -14
rect 60 -24 61 -20
rect 63 -16 68 -14
rect 63 -20 64 -16
rect 63 -24 68 -20
<< pdiffusion >>
rect 39 40 44 49
rect -9 36 -8 40
rect -13 0 -8 36
rect -6 0 2 40
rect 4 4 12 40
rect 4 0 6 4
rect 10 0 12 4
rect 14 36 15 40
rect 14 0 19 36
rect 23 4 28 40
rect 27 0 28 4
rect 30 36 31 40
rect 35 36 36 40
rect 30 0 36 36
rect 38 0 45 40
rect 60 14 61 18
rect 56 -2 61 14
rect 63 4 68 18
rect 63 0 64 4
rect 63 -2 68 0
<< metal1 >>
rect -9 56 -5 59
rect 1 56 5 59
rect 11 56 15 59
rect 27 56 31 59
rect 35 56 39 59
rect -13 40 -9 44
rect 19 36 31 40
rect 56 18 60 22
rect 6 -5 10 0
rect 23 -5 27 0
rect 64 -5 68 0
rect -4 -9 57 -5
rect 64 -9 75 -5
rect -4 -14 0 -9
rect 10 -18 39 -14
rect 64 -16 68 -9
rect 56 -28 60 -24
rect 19 -34 23 -30
rect -13 -42 -9 -34
rect 31 -38 35 -34
rect -5 -42 35 -38
<< metal2 >>
rect -5 44 44 49
rect -5 39 0 44
rect 39 39 44 44
<< ntransistor >>
rect -8 -34 -6 -14
rect 2 -34 4 -14
rect 12 -34 14 -14
rect 28 -34 30 -14
rect 36 -34 38 -14
rect 61 -24 63 -14
<< ptransistor >>
rect -8 0 -6 40
rect 2 0 4 40
rect 12 0 14 40
rect 28 0 30 40
rect 36 0 38 40
rect 61 -2 63 18
<< polycontact >>
rect -9 52 -5 56
rect 1 52 5 56
rect 11 52 15 56
rect 27 52 31 56
rect 35 52 39 56
rect 57 -9 61 -5
<< ndcontact >>
rect -13 -34 -9 -30
rect -4 -18 0 -14
rect 6 -18 10 -14
rect 15 -34 19 -30
rect 23 -34 27 -30
rect 31 -34 35 -30
rect 39 -18 43 -14
rect 56 -24 60 -20
rect 64 -20 68 -16
<< pdcontact >>
rect -13 36 -9 40
rect 6 0 10 4
rect 15 36 19 40
rect 23 0 27 4
rect 31 36 35 40
rect 56 14 60 18
rect 64 0 68 4
<< m2contact >>
rect -5 34 0 39
rect 39 34 44 39
<< psubstratepcontact >>
rect 56 -32 60 -28
rect -9 -42 -5 -38
<< nsubstratencontact >>
rect -13 44 -9 48
rect 56 22 60 26
<< labels >>
rlabel metal1 -13 -40 -11 -39 1 gnd
rlabel nsubstratencontact -12 44 -10 45 1 vdd
rlabel metal1 -8 57 -6 58 5 G2
rlabel metal1 2 57 4 58 5 P2
rlabel metal1 12 57 14 58 5 P1
rlabel metal1 28 57 30 58 5 G0
rlabel metal1 36 57 38 58 5 G1
rlabel metal1 56 20 60 21 1 vdd
rlabel metal1 56 -28 60 -27 1 gnd
rlabel metal1 49 -8 50 -6 1 C3_bar
rlabel metal1 74 -8 75 -6 7 C3
<< end >>
