* SPICE3 file created from C5.ext - technology: scmos

.option scale=90n

M1000 a_n7_0# G0 gnd Gnd nfet w=20 l=2
+  ad=80p pd=28u as=100p ps=50u
M1001 a_13_0# P2 a_3_0# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=80p ps=28u
M1002 C5_bar P4 a_49_0# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=80p ps=28u
M1003 a_49_0# P3 a_13_0# Gnd nfet w=20 l=2
+  ad=80p pd=28u as=80p ps=28u
M1004 a_13_0# G2 gnd Gnd nfet w=20 l=2
+  ad=80p pd=28u as=80p ps=28u
M1005 gnd G1 a_3_0# Gnd nfet w=20 l=2
+  ad=80p pd=28u as=100p ps=50u
M1006 C5_bar G4 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=80p ps=28u
M1007 gnd G3 a_49_0# Gnd nfet w=20 l=2
+  ad=80p pd=28u as=100p ps=50u
M1008 a_13_34# G1 a_n7_34# vdd pfet w=40 l=2
+  ad=0.16n pd=48u as=0.2n ps=90u
M1009 C5 C5_bar vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1010 C5 C5_bar gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M1011 a_13_34# P2 vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.16n ps=48u
M1012 a_59_34# G3 a_39_34# vdd pfet w=40 l=2
+  ad=0.16n pd=48u as=0.2n ps=90u
M1013 a_n7_34# G0 vdd vdd pfet w=40 l=2
+  ad=0.16n pd=48u as=0.2n ps=90u
M1014 a_39_34# G2 a_13_34# vdd pfet w=40 l=2
+  ad=0.16n pd=48u as=0.16n ps=48u
M1015 C5_bar G4 a_59_34# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.16n ps=48u
M1016 vdd P1 a_n7_34# vdd pfet w=40 l=2
+  ad=0.16n pd=48u as=0.16n ps=48u
M1017 vdd P3 a_39_34# vdd pfet w=40 l=2
+  ad=0.16n pd=48u as=0.16n ps=48u
M1018 a_3_0# P1 a_n7_0# Gnd nfet w=20 l=2
+  ad=80p pd=28u as=80p ps=28u
M1019 a_59_34# P4 vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.16n ps=48u
C0 vdd 0 8.07907f