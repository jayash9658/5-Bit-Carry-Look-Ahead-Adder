magic
tech scmos
timestamp 1763289728
<< nwell >>
rect -18 -6 13 31
<< ntransistor >>
rect -5 -22 -3 -12
<< ptransistor >>
rect -5 0 -3 20
<< ndiffusion >>
rect -10 -18 -5 -12
rect -6 -22 -5 -18
rect -3 -14 2 -12
rect -3 -18 -2 -14
rect -3 -22 2 -18
<< pdiffusion >>
rect -6 16 -5 20
rect -10 0 -5 16
rect -3 6 2 20
rect -3 2 -2 6
rect -3 0 2 2
<< ndcontact >>
rect -10 -22 -6 -18
rect -2 -18 2 -14
<< pdcontact >>
rect -10 16 -6 20
rect -2 2 2 6
<< psubstratepcontact >>
rect -10 -30 -6 -26
<< nsubstratencontact >>
rect -10 24 -6 28
<< polysilicon >>
rect -5 20 -3 23
rect -5 -12 -3 0
rect -5 -25 -3 -22
<< polycontact >>
rect -9 -7 -5 -3
<< metal1 >>
rect -10 20 -6 24
rect -2 -3 2 2
rect -17 -7 -9 -3
rect -2 -7 9 -3
rect -2 -14 2 -7
rect -10 -26 -6 -22
<< labels >>
rlabel metal1 -17 -6 -16 -4 3 Vin
rlabel metal1 8 -6 9 -4 7 Vout
rlabel metal1 -10 22 -6 23 1 vdd
rlabel metal1 -10 -26 -6 -25 1 gnd
<< end >>
