magic
tech scmos
timestamp 1763293589
<< nwell >>
rect -20 30 19 31
rect -20 -6 46 30
rect 16 -7 46 -6
<< ntransistor >>
rect -9 -22 -7 -12
rect 3 -22 5 -12
rect 28 -23 30 -13
<< ptransistor >>
rect -9 0 -7 20
rect 3 0 5 20
rect 28 -1 30 19
<< ndiffusion >>
rect -14 -18 -9 -12
rect -10 -22 -9 -18
rect -7 -22 3 -12
rect 5 -16 6 -12
rect 5 -22 10 -16
rect 23 -19 28 -13
rect 27 -23 28 -19
rect 30 -15 35 -13
rect 30 -19 31 -15
rect 30 -23 35 -19
<< pdiffusion >>
rect -10 16 -9 20
rect -14 0 -9 16
rect -7 5 3 20
rect -7 1 -4 5
rect 0 1 3 5
rect -7 0 3 1
rect 5 16 6 20
rect 5 0 10 16
rect 27 15 28 19
rect 23 -1 28 15
rect 30 5 35 19
rect 30 1 31 5
rect 30 -1 35 1
<< ndcontact >>
rect -14 -22 -10 -18
rect 6 -16 10 -12
rect 23 -23 27 -19
rect 31 -19 35 -15
<< pdcontact >>
rect -14 16 -10 20
rect -4 1 0 5
rect 6 16 10 20
rect 23 15 27 19
rect 31 1 35 5
<< psubstratepcontact >>
rect -14 -30 -10 -26
rect 23 -31 27 -27
<< nsubstratencontact >>
rect -4 24 0 28
rect 23 23 27 27
<< polysilicon >>
rect -9 20 -7 31
rect 3 20 5 31
rect 28 19 30 22
rect -9 -12 -7 0
rect 3 -12 5 0
rect 28 -13 30 -1
rect -9 -25 -7 -22
rect 3 -25 5 -22
rect 28 -26 30 -23
<< polycontact >>
rect -10 31 -6 35
rect 2 31 6 35
rect 24 -8 28 -4
<< metal1 >>
rect -10 35 -6 39
rect 2 35 6 39
rect -14 24 -4 28
rect 0 24 10 28
rect -14 20 -10 24
rect 6 20 10 24
rect 23 19 27 23
rect -4 -4 0 1
rect 31 -4 35 1
rect -4 -8 24 -4
rect 31 -8 42 -4
rect 6 -12 10 -8
rect 31 -15 35 -8
rect -14 -26 -10 -22
rect 23 -27 27 -23
<< labels >>
rlabel metal1 -14 -26 -13 -24 2 gnd
rlabel metal1 -14 27 -10 28 5 vdd
rlabel metal1 -9 38 -7 39 5 B
rlabel metal1 3 38 5 39 5 A
rlabel metal1 23 21 27 22 1 vdd
rlabel metal1 23 -27 27 -26 1 gnd
rlabel metal1 13 -7 18 -6 1 Y_bar
rlabel metal1 41 -7 42 -5 7 Y
<< end >>
