.include TSMC_180nm.txt
.include INV.sp
.param LAMBDA=0.09u
.param Width_N = 10*LAMBDA
.param Width_P = 20*LAMBDA
.global vdd gnd

Vdd vdd 0 1.8
Vclk clk 0 pulse(0 1.8 0 100p 100p 10n 20n)
Vdata D 0 pwl(0 0 12n 0 12.1n 1.8 32n 1.8 32.1n 0 60n 0)


M3 l1 D vdd vdd CMOSP W={Width_P} L={2*LAMBDA}
+ AS={5*Width_P*LAMBDA} PS={10*LAMBDA+2*Width_P}
+ AD={5*Width_P*LAMBDA} PD={10*LAMBDA+2*Width_P}
M2 X clk l1 vdd CMOSP W={Width_P} L={2*LAMBDA}
+ AS={5*Width_P*LAMBDA} PS={10*LAMBDA+2*Width_P}
+ AD={5*Width_P*LAMBDA} PD={10*LAMBDA+2*Width_P}
M1 X D gnd gnd CMOSN W={Width_N} L={2*LAMBDA}
+ AS={5*Width_N*LAMBDA} PS={10*LAMBDA+2*Width_N}
+ AD={5*Width_N*LAMBDA} PD={10*LAMBDA+2*Width_N}

M6 Y clk vdd vdd CMOSP W={Width_P} L={2*LAMBDA}
+ AS={5*Width_P*LAMBDA} PS={10*LAMBDA+2*Width_P}
+ AD={5*Width_P*LAMBDA} PD={10*LAMBDA+2*Width_P}
M5 Y X l2 gnd CMOSN W={Width_N} L={2*LAMBDA}
+ AS={5*Width_N*LAMBDA} PS={10*LAMBDA+2*Width_N}
+ AD={5*Width_N*LAMBDA} PD={10*LAMBDA+2*Width_N}
M4 l2 clk gnd gnd CMOSN W={Width_N} L={2*LAMBDA}
+ AS={5*Width_N*LAMBDA} PS={10*LAMBDA+2*Width_N}
+ AD={5*Width_N*LAMBDA} PD={10*LAMBDA+2*Width_N}

M9 Q_bar Y vdd vdd CMOSP W={Width_P} L={2*LAMBDA}
+ AS={5*Width_P*LAMBDA} PS={10*LAMBDA+2*Width_P}
+ AD={5*Width_P*LAMBDA} PD={10*LAMBDA+2*Width_P}
M8 Q_bar clk l3 gnd CMOSN W={Width_N} L={2*LAMBDA}
+ AS={5*Width_N*LAMBDA} PS={10*LAMBDA+2*Width_N}
+ AD={5*Width_N*LAMBDA} PD={10*LAMBDA+2*Width_N}
M7 l3 Y gnd gnd CMOSN W={Width_N} L={2*LAMBDA}
+ AS={5*Width_N*LAMBDA} PS={10*LAMBDA+2*Width_N}
+ AD={5*Width_N*LAMBDA} PD={10*LAMBDA+2*Width_N}

x1 Q Q_bar vdd gnd inv


.tran 0.01n 60n
.measure tran tcpq
+ TRIG v(clk) VAL=0.9 RISE=2
+ TARG v(Q) VAL=0.9 RISE=1

.measure tran tsetup
+ TRIG v(D) VAL=0.9 RISE=1
+ TARG v(X) VAL=0.9 FALL=1

.measure tran thold
+ TRIG v(Y) VAL=0.9 FALL=1
+ TARG v(X) VAL=0.9 RISE=1

.control
run
plot clk D+2 Q+4 X+6 Y+8
.endc

.end