magic
tech scmos
timestamp 1764588473
<< checkpaint >>
rect 170760400 14000 869359811 25949
rect 170760800 400 869359811 14000
rect 54 143 869359811 400
rect -16 138 869359811 143
rect -63 135 869359811 138
rect -70 134 869359811 135
rect -104 -7 869359811 134
rect -104 -9 477026675 -7
rect -104 -67 226 -9
rect 30196400 -67 477026675 -9
rect -104 -70 148 -67
rect -57 -75 89 -70
<< nwell >>
rect 32 357 80 378
rect 23 300 80 357
rect 206 333 243 364
rect 38 276 80 300
rect 179 330 243 333
rect 179 286 244 330
rect 327 272 375 293
rect 9 238 46 265
rect 8 235 46 238
rect 8 199 45 235
rect 318 215 375 272
rect 333 191 375 215
rect 32 158 80 179
rect 23 101 80 158
rect 38 77 80 101
rect 8 39 45 66
rect 7 36 45 39
rect 7 3 44 36
rect 14 0 44 3
<< ntransistor >>
rect 88 360 98 362
rect 249 346 259 348
rect 86 344 106 346
rect 86 336 106 338
rect 86 328 106 330
rect 86 319 106 321
rect 252 317 272 319
rect 252 307 272 309
rect 88 295 98 297
rect 252 297 272 299
rect 383 275 393 277
rect 381 259 401 261
rect 381 251 401 253
rect 52 247 62 249
rect 381 243 401 245
rect 381 234 401 236
rect 51 222 61 224
rect 51 210 61 212
rect 383 210 393 212
rect 88 161 98 163
rect 86 145 106 147
rect 86 137 106 139
rect 86 129 106 131
rect 86 120 106 122
rect 88 96 98 98
rect 51 48 61 50
rect 50 23 60 25
rect 50 11 60 13
<< ptransistor >>
rect 49 360 69 362
rect 217 346 237 348
rect 29 344 69 346
rect 29 336 69 338
rect 29 328 69 330
rect 29 319 69 321
rect 198 317 238 319
rect 198 307 238 309
rect 49 295 69 297
rect 198 297 238 299
rect 344 275 364 277
rect 324 259 364 261
rect 324 251 364 253
rect 20 247 40 249
rect 324 243 364 245
rect 324 234 364 236
rect 19 222 39 224
rect 19 210 39 212
rect 344 210 364 212
rect 49 161 69 163
rect 29 145 69 147
rect 29 137 69 139
rect 29 129 69 131
rect 29 120 69 122
rect 49 96 69 98
rect 19 48 39 50
rect 18 23 38 25
rect 18 11 38 13
<< ndiffusion >>
rect 88 364 90 368
rect 94 364 98 368
rect 88 362 98 364
rect 88 359 98 360
rect 88 355 94 359
rect 90 347 106 351
rect 249 349 251 353
rect 255 349 259 353
rect 249 348 259 349
rect 86 346 106 347
rect 86 338 106 344
rect 249 345 259 346
rect 249 341 255 345
rect 86 335 106 336
rect 86 331 102 335
rect 86 330 106 331
rect 86 321 106 328
rect 86 318 106 319
rect 90 314 106 318
rect 252 320 268 324
rect 252 319 272 320
rect 252 315 272 317
rect 256 311 272 315
rect 252 309 272 311
rect 92 298 98 302
rect 88 297 98 298
rect 252 299 272 307
rect 88 293 98 295
rect 88 289 94 293
rect 252 296 272 297
rect 252 292 268 296
rect 383 279 385 283
rect 389 279 393 283
rect 383 277 393 279
rect 383 274 393 275
rect 383 270 389 274
rect 385 262 401 266
rect 381 261 401 262
rect 52 250 54 254
rect 58 250 62 254
rect 381 253 401 259
rect 52 249 62 250
rect 52 246 62 247
rect 52 242 58 246
rect 381 250 401 251
rect 381 246 397 250
rect 381 245 401 246
rect 381 236 401 243
rect 381 233 401 234
rect 385 229 401 233
rect 55 225 61 229
rect 51 224 61 225
rect 51 212 61 222
rect 51 209 61 210
rect 387 213 393 217
rect 383 212 393 213
rect 51 205 57 209
rect 383 208 393 210
rect 383 204 389 208
rect 88 165 90 169
rect 94 165 98 169
rect 88 163 98 165
rect 88 160 98 161
rect 88 156 94 160
rect 90 148 106 152
rect 86 147 106 148
rect 86 139 106 145
rect 86 136 106 137
rect 86 132 102 136
rect 86 131 106 132
rect 86 122 106 129
rect 86 119 106 120
rect 90 115 106 119
rect 92 99 98 103
rect 88 98 98 99
rect 88 94 98 96
rect 88 90 94 94
rect 51 51 53 55
rect 57 51 61 55
rect 51 50 61 51
rect 51 47 61 48
rect 51 43 57 47
rect 54 26 60 30
rect 50 25 60 26
rect 50 13 60 23
rect 50 10 60 11
rect 50 6 56 10
<< pdiffusion >>
rect 49 364 63 368
rect 67 364 69 368
rect 49 362 69 364
rect 49 359 69 360
rect 49 355 65 359
rect 49 354 69 355
rect 33 347 69 351
rect 29 346 69 347
rect 217 349 231 353
rect 235 349 237 353
rect 217 348 237 349
rect 217 345 237 346
rect 29 343 69 344
rect 29 339 65 343
rect 29 338 69 339
rect 221 341 237 345
rect 29 335 69 336
rect 33 331 69 335
rect 29 330 69 331
rect 29 326 69 328
rect 29 322 65 326
rect 29 321 69 322
rect 198 320 234 324
rect 29 318 69 319
rect 33 314 69 318
rect 198 319 238 320
rect 198 315 238 317
rect 198 311 234 315
rect 198 309 238 311
rect 198 305 238 307
rect 49 302 69 303
rect 49 298 65 302
rect 49 297 69 298
rect 202 301 238 305
rect 198 299 238 301
rect 198 296 238 297
rect 49 293 69 295
rect 49 289 65 293
rect 198 292 234 296
rect 344 279 358 283
rect 362 279 364 283
rect 344 277 364 279
rect 344 274 364 275
rect 344 270 360 274
rect 344 269 364 270
rect 328 262 364 266
rect 324 261 364 262
rect 324 258 364 259
rect 324 254 360 258
rect 20 250 34 254
rect 38 250 40 254
rect 20 249 40 250
rect 324 253 364 254
rect 324 250 364 251
rect 20 246 40 247
rect 24 242 40 246
rect 328 246 364 250
rect 324 245 364 246
rect 324 241 364 243
rect 324 237 360 241
rect 324 236 364 237
rect 324 233 364 234
rect 328 229 364 233
rect 23 225 39 229
rect 19 224 39 225
rect 19 219 39 222
rect 19 215 34 219
rect 38 215 39 219
rect 19 212 39 215
rect 344 217 364 218
rect 344 213 360 217
rect 19 209 39 210
rect 23 205 39 209
rect 344 212 364 213
rect 344 208 364 210
rect 344 204 360 208
rect 49 165 63 169
rect 67 165 69 169
rect 49 163 69 165
rect 49 160 69 161
rect 49 156 65 160
rect 49 155 69 156
rect 33 148 69 152
rect 29 147 69 148
rect 29 144 69 145
rect 29 140 65 144
rect 29 139 69 140
rect 29 136 69 137
rect 33 132 69 136
rect 29 131 69 132
rect 29 127 69 129
rect 29 123 65 127
rect 29 122 69 123
rect 29 119 69 120
rect 33 115 69 119
rect 49 103 69 104
rect 49 99 65 103
rect 49 98 69 99
rect 49 94 69 96
rect 49 90 65 94
rect 19 51 33 55
rect 37 51 39 55
rect 19 50 39 51
rect 19 47 39 48
rect 23 43 39 47
rect 22 26 38 30
rect 18 25 38 26
rect 18 20 38 23
rect 18 16 33 20
rect 37 16 38 20
rect 18 13 38 16
rect 18 10 38 11
rect 22 6 38 10
<< ndcontact >>
rect 90 364 94 368
rect 94 355 98 359
rect 86 347 90 351
rect 251 349 255 353
rect 255 341 259 345
rect 102 331 106 335
rect 86 314 90 318
rect 268 320 272 324
rect 252 311 256 315
rect 88 298 92 302
rect 94 289 98 293
rect 268 292 272 296
rect 385 279 389 283
rect 389 270 393 274
rect 381 262 385 266
rect 54 250 58 254
rect 58 242 62 246
rect 397 246 401 250
rect 381 229 385 233
rect 51 225 55 229
rect 383 213 387 217
rect 57 205 61 209
rect 389 204 393 208
rect 90 165 94 169
rect 94 156 98 160
rect 86 148 90 152
rect 102 132 106 136
rect 86 115 90 119
rect 88 99 92 103
rect 94 90 98 94
rect 53 51 57 55
rect 57 43 61 47
rect 50 26 54 30
rect 56 6 60 10
<< pdcontact >>
rect 63 364 67 368
rect 65 355 69 359
rect 29 347 33 351
rect 231 349 235 353
rect 65 339 69 343
rect 217 341 221 345
rect 29 331 33 335
rect 123 331 127 335
rect 65 322 69 326
rect 234 320 238 324
rect 29 314 33 318
rect 234 311 238 315
rect 65 298 69 302
rect 198 301 202 305
rect 65 289 69 293
rect 234 292 238 296
rect 358 279 362 283
rect 360 270 364 274
rect 324 262 328 266
rect 360 254 364 258
rect 34 250 38 254
rect 20 242 24 246
rect 324 246 328 250
rect 418 246 422 250
rect 360 237 364 241
rect 324 229 328 233
rect 19 225 23 229
rect 34 215 38 219
rect 360 213 364 217
rect 19 205 23 209
rect 360 204 364 208
rect 63 165 67 169
rect 65 156 69 160
rect 29 148 33 152
rect 65 140 69 144
rect 29 132 33 136
rect 123 132 127 136
rect 65 123 69 127
rect 29 115 33 119
rect 65 99 69 103
rect 65 90 69 94
rect 33 51 37 55
rect 19 43 23 47
rect 18 26 22 30
rect 33 16 37 20
rect 18 6 22 10
<< psubstratepcontact >>
rect 263 341 267 345
rect 110 331 114 335
rect 276 301 280 305
rect 66 242 70 246
rect 405 246 409 250
rect 65 205 69 209
rect 110 132 114 136
rect 65 43 69 47
rect 64 6 68 10
<< nsubstratencontact >>
rect 209 341 213 345
rect 190 301 194 305
rect 65 279 69 283
rect 12 242 16 246
rect 11 215 15 219
rect 360 194 364 198
rect 65 80 69 84
rect 11 43 15 47
rect 10 16 14 20
<< polysilicon >>
rect 48 360 49 362
rect 69 360 88 362
rect 98 360 101 362
rect 214 346 217 348
rect 237 346 249 348
rect 259 346 262 348
rect 1 344 29 346
rect 69 344 86 346
rect 106 344 109 346
rect 17 336 29 338
rect 69 336 86 338
rect 106 336 109 338
rect 0 328 29 330
rect 69 328 86 330
rect 106 328 109 330
rect 1 319 29 321
rect 69 319 86 321
rect 106 319 109 321
rect 187 317 198 319
rect 238 317 252 319
rect 272 317 275 319
rect 187 307 198 309
rect 238 307 252 309
rect 272 307 275 309
rect 48 295 49 297
rect 69 295 88 297
rect 98 295 101 297
rect 187 297 198 299
rect 238 297 252 299
rect 272 297 275 299
rect 343 275 344 277
rect 364 275 383 277
rect 393 275 396 277
rect 296 259 324 261
rect 364 259 381 261
rect 401 259 404 261
rect 312 251 324 253
rect 364 251 381 253
rect 401 251 404 253
rect 17 247 20 249
rect 40 247 52 249
rect 62 247 65 249
rect 295 243 324 245
rect 364 243 381 245
rect 401 243 404 245
rect 296 234 324 236
rect 364 234 381 236
rect 401 234 404 236
rect 8 222 19 224
rect 39 222 51 224
rect 61 222 64 224
rect 8 210 19 212
rect 39 210 51 212
rect 61 210 64 212
rect 343 210 344 212
rect 364 210 383 212
rect 393 210 396 212
rect 48 161 49 163
rect 69 161 88 163
rect 98 161 101 163
rect 1 145 29 147
rect 69 145 86 147
rect 106 145 109 147
rect 17 137 29 139
rect 69 137 86 139
rect 106 137 109 139
rect 0 129 29 131
rect 69 129 86 131
rect 106 129 109 131
rect 1 120 29 122
rect 69 120 86 122
rect 106 120 109 122
rect 48 96 49 98
rect 69 96 88 98
rect 98 96 101 98
rect 16 48 19 50
rect 39 48 51 50
rect 61 48 64 50
rect 7 23 18 25
rect 38 23 50 25
rect 60 23 63 25
rect 7 11 18 13
rect 38 11 50 13
rect 60 11 63 13
<< polycontact >>
rect 44 359 48 363
rect -3 343 1 347
rect 13 335 17 339
rect 240 342 244 346
rect -4 327 0 331
rect -3 318 1 322
rect 183 316 187 320
rect 183 306 187 310
rect 44 294 48 298
rect 183 296 187 300
rect 339 274 343 278
rect 292 258 296 262
rect 308 250 312 254
rect 43 243 47 247
rect 291 242 295 246
rect 292 233 296 237
rect 4 221 8 225
rect 4 209 8 213
rect 339 209 343 213
rect 44 160 48 164
rect -3 144 1 148
rect 13 136 17 140
rect -4 128 0 132
rect -3 119 1 123
rect 44 95 48 99
rect 42 44 46 48
rect 3 22 7 26
rect 3 10 7 14
<< metal1 >>
rect -3 371 76 375
rect -3 347 1 371
rect 72 368 76 371
rect 67 364 90 368
rect 5 359 44 363
rect -4 331 0 334
rect 5 322 9 359
rect 69 355 72 359
rect 98 355 114 359
rect 21 347 29 351
rect 1 318 9 322
rect 13 310 17 335
rect 21 335 25 347
rect 81 343 85 347
rect 69 339 85 343
rect 21 331 29 335
rect 21 318 25 331
rect 69 322 72 326
rect 81 318 85 339
rect 110 335 114 355
rect 240 353 244 360
rect 235 349 251 353
rect 213 341 217 345
rect 106 331 110 335
rect 114 331 123 335
rect 21 314 29 318
rect 81 314 86 318
rect 13 306 84 310
rect 80 302 84 306
rect 69 298 88 302
rect 9 294 44 298
rect 69 289 72 293
rect 110 293 114 331
rect 240 324 244 342
rect 259 341 263 345
rect 238 320 251 324
rect 272 320 280 324
rect 98 289 114 293
rect 165 316 183 320
rect 65 283 69 289
rect 165 261 169 316
rect 247 315 251 320
rect 238 311 243 315
rect 247 311 252 315
rect 181 306 183 310
rect 194 301 198 305
rect 43 257 169 261
rect 172 296 183 300
rect 239 296 243 311
rect 276 305 280 320
rect 276 296 280 301
rect 43 254 47 257
rect 38 250 54 254
rect 16 242 20 246
rect 43 229 47 243
rect 62 242 66 246
rect 172 237 176 296
rect 238 292 243 296
rect 272 292 280 296
rect 292 286 371 290
rect 292 262 296 286
rect 367 283 371 286
rect 362 279 385 283
rect 300 274 339 278
rect 291 246 295 249
rect 300 237 304 274
rect 364 270 367 274
rect 393 270 409 274
rect 316 262 324 266
rect 172 233 292 237
rect 296 233 304 237
rect 308 237 312 250
rect 316 250 320 262
rect 376 258 380 262
rect 364 254 380 258
rect 316 246 324 250
rect 316 237 320 246
rect 364 237 367 241
rect 308 233 314 237
rect 316 233 322 237
rect 376 233 380 254
rect 405 250 409 270
rect 401 246 405 250
rect 409 246 418 250
rect 11 225 19 229
rect 43 225 51 229
rect 0 221 4 225
rect 11 219 15 225
rect 43 219 47 225
rect 38 215 47 219
rect 0 209 4 213
rect 11 209 15 215
rect 11 205 19 209
rect 61 205 65 209
rect -3 172 76 176
rect -3 148 1 172
rect 72 169 76 172
rect 67 165 90 169
rect 5 160 44 164
rect -4 132 0 135
rect 5 123 9 160
rect 69 156 72 160
rect 98 156 114 160
rect 21 148 29 152
rect 1 119 9 123
rect 13 111 17 136
rect 21 136 25 148
rect 81 144 85 148
rect 69 140 85 144
rect 21 132 29 136
rect 21 119 25 132
rect 69 123 72 127
rect 81 119 85 140
rect 110 136 114 156
rect 106 132 110 136
rect 114 132 123 136
rect 21 115 29 119
rect 81 115 86 119
rect 13 107 84 111
rect 80 103 84 107
rect 69 99 88 103
rect 9 95 44 99
rect 69 90 72 94
rect 110 94 114 132
rect 98 90 114 94
rect 65 84 69 90
rect 172 62 176 233
rect 308 225 312 233
rect 316 229 324 233
rect 376 229 381 233
rect 308 221 379 225
rect 375 217 379 221
rect 364 213 383 217
rect 304 209 339 213
rect 364 204 367 208
rect 405 208 409 246
rect 393 204 409 208
rect 360 198 364 204
rect 42 58 176 62
rect 42 55 46 58
rect 37 51 53 55
rect 15 43 19 47
rect 42 30 46 44
rect 61 43 65 47
rect 10 26 18 30
rect 42 26 50 30
rect -1 22 3 26
rect 10 20 14 26
rect 42 20 46 26
rect 37 16 46 20
rect -1 10 3 14
rect 10 10 14 16
rect 10 6 18 10
rect 60 6 64 10
<< m2contact >>
rect -5 334 0 339
rect 72 354 77 359
rect 81 347 86 352
rect 72 322 77 327
rect 4 294 9 299
rect 72 289 77 294
rect 176 306 181 311
rect 290 249 295 254
rect 367 269 372 274
rect 376 262 381 267
rect 367 237 372 242
rect -5 135 0 140
rect 72 155 77 160
rect 81 148 86 153
rect 72 123 77 128
rect 4 95 9 100
rect 72 90 77 95
rect 299 209 304 214
rect 367 204 372 209
<< metal2 >>
rect 81 370 162 375
rect 0 335 9 339
rect 4 299 9 335
rect 73 327 77 354
rect 81 352 86 370
rect 73 294 77 322
rect 157 311 162 370
rect 157 306 176 311
rect 157 254 162 306
rect 376 292 450 297
rect 157 249 290 254
rect 295 250 304 254
rect 299 249 305 250
rect 310 249 322 254
rect 299 214 304 249
rect 368 242 372 269
rect 376 267 381 292
rect 368 209 372 237
rect 81 175 419 180
rect 0 136 9 140
rect 4 100 9 136
rect 73 128 77 155
rect 81 153 86 175
rect 73 95 77 123
<< labels >>
rlabel metal1 108 132 114 136 7 gnd
rlabel metal1 101 156 102 160 7 gnd
rlabel nsubstratencontact 65 80 69 84 1 vdd
rlabel metal1 63 205 65 206 8 gnd
rlabel metal1 11 205 12 209 3 vdd
rlabel metal1 17 242 18 246 7 vdd
rlabel metal1 65 242 66 246 7 gnd
rlabel metal1 108 331 114 335 7 gnd
rlabel metal1 101 355 102 359 7 gnd
rlabel nsubstratencontact 65 279 69 283 1 vdd
rlabel polycontact -3 119 1 123 3 A0
rlabel polycontact -4 128 0 132 3 B0
rlabel metal1 0 210 1 212 3 B1
rlabel metal1 0 222 1 224 3 A1
rlabel polycontact -3 318 1 322 3 A1
rlabel polycontact -4 327 0 331 3 B1
rlabel metal1 190 301 191 304 3 vdd
rlabel metal1 181 296 182 299 3 G0
rlabel metal1 181 316 182 319 3 G1
rlabel metal1 214 341 215 345 7 vdd
rlabel metal1 262 341 263 345 7 gnd
rlabel metal1 242 328 243 333 7 C2_bar
rlabel metal1 241 359 243 360 5 C2
rlabel metal1 277 292 278 295 8 gnd
rlabel metal1 181 306 182 309 3 P1
rlabel metal2 445 292 450 297 7 S1
rlabel metal2 414 175 419 180 1 S0
rlabel nsubstratencontact 360 194 364 198 1 vdd
rlabel metal1 396 270 397 274 7 gnd
rlabel metal1 403 246 409 250 7 gnd
rlabel polycontact 13 136 17 140 1 B0_bar
rlabel polycontact -3 144 1 148 3 A0_bar
rlabel metal1 45 232 46 237 1 G1_bar
rlabel polycontact 13 335 17 339 1 B1_bar
rlabel polycontact -3 343 1 347 3 A1_bar
rlabel polycontact 291 242 295 246 1 P1
rlabel polycontact 292 233 296 237 1 G0
rlabel polycontact 292 258 296 262 1 G0_bar
rlabel polycontact 308 250 312 254 1 P1_bar
rlabel metal1 62 6 64 7 8 gnd
rlabel metal1 10 6 11 10 3 vdd
rlabel metal1 16 43 17 47 7 vdd
rlabel metal1 64 43 65 47 7 gnd
rlabel metal1 44 33 45 38 1 G0_bar
rlabel metal1 -1 11 0 13 3 B0
rlabel metal1 -1 23 0 25 3 A0
<< end >>
