magic
tech scmos
timestamp 1764625264
<< checkpaint >>
rect 579159200 5200 869359811 25949
rect 579159600 400 869359811 5200
rect -183 -7 869359811 400
rect -183 -9 477026675 -7
rect -567 -193 -430 -56
rect -183 -99 905 -9
rect 1289 -84 1550 -9
rect 30196400 -67 477026675 -9
rect -183 -132 23 -99
rect 40 -108 402 -99
rect 40 -110 279 -108
rect 40 -175 249 -110
rect 40 -310 178 -175
<< nwell >>
rect -8 948 40 969
rect -17 891 40 948
rect 241 920 278 951
rect -2 872 40 891
rect 18 867 40 872
rect -35 828 2 855
rect -36 825 2 828
rect -36 789 1 825
rect 217 804 275 920
rect 374 815 422 836
rect -8 753 40 774
rect 365 758 422 815
rect -17 696 40 753
rect 241 710 278 741
rect 380 734 422 758
rect -2 677 40 696
rect 18 672 40 677
rect -35 628 2 655
rect -36 625 2 628
rect -36 589 1 625
rect 217 614 275 710
rect 374 621 422 642
rect -8 555 40 576
rect 365 564 422 621
rect -17 498 40 555
rect 380 540 422 564
rect -2 479 40 498
rect 18 474 40 479
rect 216 489 279 520
rect -35 434 2 461
rect -36 431 2 434
rect -36 395 1 431
rect 216 422 278 489
rect 374 408 422 429
rect -8 357 40 378
rect -17 300 40 357
rect 365 351 422 408
rect 380 327 422 351
rect -2 276 40 300
rect 242 284 279 315
rect 215 281 279 284
rect -35 237 2 264
rect 215 237 280 281
rect 374 254 422 275
rect -36 234 2 237
rect -36 198 1 234
rect 365 197 422 254
rect -8 154 40 175
rect 380 173 422 197
rect -17 97 40 154
rect -2 78 40 97
rect 18 73 40 78
rect -35 22 2 49
rect -36 19 2 22
rect -36 -17 1 19
<< ntransistor >>
rect 48 951 58 953
rect 46 935 66 937
rect 284 933 294 935
rect 46 927 66 929
rect 46 919 66 921
rect 46 910 66 912
rect 283 907 303 909
rect 283 897 303 899
rect 48 886 58 888
rect 283 881 303 883
rect 283 871 303 873
rect 283 861 303 863
rect 283 851 303 853
rect 8 837 18 839
rect 283 835 303 837
rect 283 825 303 827
rect 430 818 440 820
rect 283 815 303 817
rect 7 812 17 814
rect 7 800 17 802
rect 428 802 448 804
rect 428 794 448 796
rect 428 786 448 788
rect 428 777 448 779
rect 48 756 58 758
rect 430 753 440 755
rect 46 740 66 742
rect 46 732 66 734
rect 46 724 66 726
rect 284 723 294 725
rect 46 715 66 717
rect 283 697 303 699
rect 48 691 58 693
rect 283 687 303 689
rect 283 677 303 679
rect 283 661 303 663
rect 283 651 303 653
rect 8 637 18 639
rect 283 635 303 637
rect 283 625 303 627
rect 430 624 440 626
rect 7 612 17 614
rect 428 608 448 610
rect 7 600 17 602
rect 428 600 448 602
rect 428 592 448 594
rect 428 583 448 585
rect 48 558 58 560
rect 430 559 440 561
rect 46 542 66 544
rect 46 534 66 536
rect 46 526 66 528
rect 46 517 66 519
rect 285 502 295 504
rect 48 493 58 495
rect 285 477 305 479
rect 285 469 305 471
rect 285 453 305 455
rect 8 443 18 445
rect 285 443 305 445
rect 285 433 305 435
rect 7 418 17 420
rect 430 411 440 413
rect 7 406 17 408
rect 428 395 448 397
rect 428 387 448 389
rect 428 379 448 381
rect 428 370 448 372
rect 48 360 58 362
rect 46 344 66 346
rect 430 346 440 348
rect 46 336 66 338
rect 46 328 66 330
rect 46 319 66 321
rect 285 297 295 299
rect 48 295 58 297
rect 288 268 308 270
rect 288 258 308 260
rect 8 246 18 248
rect 430 257 440 259
rect 288 248 308 250
rect 428 241 448 243
rect 428 233 448 235
rect 428 225 448 227
rect 7 221 17 223
rect 428 216 448 218
rect 7 209 17 211
rect 430 192 440 194
rect 48 157 58 159
rect 46 141 66 143
rect 46 133 66 135
rect 46 125 66 127
rect 46 116 66 118
rect 48 92 58 94
rect 8 31 18 33
rect 7 6 17 8
rect 7 -6 17 -4
<< ptransistor >>
rect 9 951 29 953
rect -11 935 29 937
rect 252 933 272 935
rect -11 927 29 929
rect -11 919 29 921
rect -11 910 29 912
rect 229 907 269 909
rect 229 897 269 899
rect 9 886 29 888
rect 229 881 269 883
rect 229 871 269 873
rect 229 861 269 863
rect 229 851 269 853
rect -24 837 -4 839
rect 229 835 269 837
rect 229 825 269 827
rect 391 818 411 820
rect 229 815 269 817
rect -25 812 -5 814
rect -25 800 -5 802
rect 371 802 411 804
rect 371 794 411 796
rect 371 786 411 788
rect 371 777 411 779
rect 9 756 29 758
rect 391 753 411 755
rect -11 740 29 742
rect -11 732 29 734
rect -11 724 29 726
rect 252 723 272 725
rect -11 715 29 717
rect 229 697 269 699
rect 9 691 29 693
rect 229 687 269 689
rect 229 677 269 679
rect 229 661 269 663
rect 229 651 269 653
rect -24 637 -4 639
rect 229 635 269 637
rect 229 625 269 627
rect 391 624 411 626
rect -25 612 -5 614
rect 371 608 411 610
rect -25 600 -5 602
rect 371 600 411 602
rect 371 592 411 594
rect 371 583 411 585
rect 9 558 29 560
rect 391 559 411 561
rect -11 542 29 544
rect -11 534 29 536
rect -11 526 29 528
rect -11 517 29 519
rect 253 502 273 504
rect 9 493 29 495
rect 231 477 271 479
rect 231 469 271 471
rect 231 453 271 455
rect -24 443 -4 445
rect 231 443 271 445
rect 231 433 271 435
rect -25 418 -5 420
rect 391 411 411 413
rect -25 406 -5 408
rect 371 395 411 397
rect 371 387 411 389
rect 371 379 411 381
rect 371 370 411 372
rect 9 360 29 362
rect -11 344 29 346
rect 391 346 411 348
rect -11 336 29 338
rect -11 328 29 330
rect -11 319 29 321
rect 253 297 273 299
rect 9 295 29 297
rect 234 268 274 270
rect 234 258 274 260
rect -24 246 -4 248
rect 391 257 411 259
rect 234 248 274 250
rect 371 241 411 243
rect 371 233 411 235
rect 371 225 411 227
rect -25 221 -5 223
rect 371 216 411 218
rect -25 209 -5 211
rect 391 192 411 194
rect 9 157 29 159
rect -11 141 29 143
rect -11 133 29 135
rect -11 125 29 127
rect -11 116 29 118
rect 9 92 29 94
rect -24 31 -4 33
rect -25 6 -5 8
rect -25 -6 -5 -4
<< ndiffusion >>
rect 48 955 50 959
rect 54 955 58 959
rect 48 953 58 955
rect 48 950 58 951
rect 48 946 54 950
rect 50 938 66 942
rect 46 937 66 938
rect 284 936 286 940
rect 290 936 294 940
rect 284 935 294 936
rect 46 929 66 935
rect 284 932 294 933
rect 284 928 290 932
rect 46 926 66 927
rect 46 922 62 926
rect 46 921 66 922
rect 46 912 66 919
rect 46 909 66 910
rect 50 905 66 909
rect 287 910 303 914
rect 283 909 303 910
rect 283 905 303 907
rect 283 901 299 905
rect 283 899 303 901
rect 52 889 58 893
rect 283 896 303 897
rect 283 892 299 896
rect 48 888 58 889
rect 48 884 58 886
rect 48 880 54 884
rect 287 884 303 888
rect 283 883 303 884
rect 283 879 303 881
rect 283 875 299 879
rect 283 873 303 875
rect 283 869 303 871
rect 287 865 303 869
rect 283 863 303 865
rect 283 859 303 861
rect 283 855 299 859
rect 283 853 303 855
rect 283 850 303 851
rect 283 846 299 850
rect 8 840 10 844
rect 14 840 18 844
rect 8 839 18 840
rect 8 836 18 837
rect 8 832 14 836
rect 287 838 303 842
rect 283 837 303 838
rect 283 833 303 835
rect 283 829 299 833
rect 283 827 303 829
rect 11 815 17 819
rect 7 814 17 815
rect 283 817 303 825
rect 430 822 432 826
rect 436 822 440 826
rect 430 820 440 822
rect 7 802 17 812
rect 283 814 303 815
rect 283 810 299 814
rect 430 817 440 818
rect 430 813 436 817
rect 432 805 448 809
rect 428 804 448 805
rect 7 799 17 800
rect 7 795 13 799
rect 428 796 448 802
rect 428 793 448 794
rect 428 789 444 793
rect 428 788 448 789
rect 428 779 448 786
rect 428 776 448 777
rect 432 772 448 776
rect 48 760 50 764
rect 54 760 58 764
rect 48 758 58 760
rect 48 755 58 756
rect 48 751 54 755
rect 434 756 440 760
rect 430 755 440 756
rect 430 751 440 753
rect 430 747 436 751
rect 50 743 66 747
rect 46 742 66 743
rect 46 734 66 740
rect 46 731 66 732
rect 46 727 62 731
rect 46 726 66 727
rect 284 726 286 730
rect 290 726 294 730
rect 284 725 294 726
rect 46 717 66 724
rect 284 722 294 723
rect 284 718 290 722
rect 46 714 66 715
rect 50 710 66 714
rect 52 694 58 698
rect 287 700 303 704
rect 283 699 303 700
rect 48 693 58 694
rect 48 689 58 691
rect 48 685 54 689
rect 283 695 303 697
rect 283 691 299 695
rect 283 689 303 691
rect 283 679 303 687
rect 283 676 303 677
rect 287 672 303 676
rect 287 664 303 668
rect 283 663 303 664
rect 283 659 303 661
rect 287 655 303 659
rect 283 653 303 655
rect 283 650 303 651
rect 283 646 299 650
rect 8 640 10 644
rect 14 640 18 644
rect 8 639 18 640
rect 8 636 18 637
rect 8 632 14 636
rect 287 638 303 642
rect 283 637 303 638
rect 283 633 303 635
rect 287 629 303 633
rect 283 627 303 629
rect 283 624 303 625
rect 283 620 299 624
rect 430 628 432 632
rect 436 628 440 632
rect 430 626 440 628
rect 430 623 440 624
rect 430 619 436 623
rect 11 615 17 619
rect 7 614 17 615
rect 7 602 17 612
rect 432 611 448 615
rect 428 610 448 611
rect 7 599 17 600
rect 428 602 448 608
rect 7 595 13 599
rect 428 599 448 600
rect 428 595 444 599
rect 428 594 448 595
rect 428 585 448 592
rect 428 582 448 583
rect 432 578 448 582
rect 48 562 50 566
rect 54 562 58 566
rect 48 560 58 562
rect 434 562 440 566
rect 430 561 440 562
rect 48 557 58 558
rect 48 553 54 557
rect 430 557 440 559
rect 430 553 436 557
rect 50 545 66 549
rect 46 544 66 545
rect 46 536 66 542
rect 46 533 66 534
rect 46 529 62 533
rect 46 528 66 529
rect 46 519 66 526
rect 46 516 66 517
rect 50 512 66 516
rect 285 505 287 509
rect 291 505 295 509
rect 285 504 295 505
rect 52 496 58 500
rect 285 501 295 502
rect 285 497 291 501
rect 48 495 58 496
rect 48 491 58 493
rect 48 487 54 491
rect 289 480 305 484
rect 285 479 305 480
rect 285 476 305 477
rect 285 472 301 476
rect 285 471 305 472
rect 285 468 305 469
rect 285 464 301 468
rect 285 456 301 460
rect 285 455 305 456
rect 8 446 10 450
rect 14 446 18 450
rect 8 445 18 446
rect 8 442 18 443
rect 285 451 305 453
rect 289 447 305 451
rect 285 445 305 447
rect 8 438 14 442
rect 285 441 305 443
rect 289 437 305 441
rect 285 435 305 437
rect 285 432 305 433
rect 285 428 301 432
rect 11 421 17 425
rect 7 420 17 421
rect 7 408 17 418
rect 430 415 432 419
rect 436 415 440 419
rect 430 413 440 415
rect 430 410 440 411
rect 430 406 436 410
rect 7 405 17 406
rect 7 401 13 405
rect 432 398 448 402
rect 428 397 448 398
rect 428 389 448 395
rect 428 386 448 387
rect 428 382 444 386
rect 428 381 448 382
rect 428 372 448 379
rect 48 364 50 368
rect 54 364 58 368
rect 428 369 448 370
rect 432 365 448 369
rect 48 362 58 364
rect 48 359 58 360
rect 48 355 54 359
rect 50 347 66 351
rect 46 346 66 347
rect 434 349 440 353
rect 430 348 440 349
rect 46 338 66 344
rect 430 344 440 346
rect 430 340 436 344
rect 46 335 66 336
rect 46 331 62 335
rect 46 330 66 331
rect 46 321 66 328
rect 46 318 66 319
rect 50 314 66 318
rect 52 298 58 302
rect 285 300 287 304
rect 291 300 295 304
rect 285 299 295 300
rect 48 297 58 298
rect 48 293 58 295
rect 48 289 54 293
rect 285 296 295 297
rect 285 292 291 296
rect 288 271 304 275
rect 288 270 308 271
rect 288 266 308 268
rect 292 262 308 266
rect 288 260 308 262
rect 8 249 10 253
rect 14 249 18 253
rect 8 248 18 249
rect 288 250 308 258
rect 430 261 432 265
rect 436 261 440 265
rect 430 259 440 261
rect 430 256 440 257
rect 430 252 436 256
rect 8 245 18 246
rect 8 241 14 245
rect 288 247 308 248
rect 288 243 304 247
rect 432 244 448 248
rect 428 243 448 244
rect 428 235 448 241
rect 11 224 17 228
rect 428 232 448 233
rect 428 228 444 232
rect 428 227 448 228
rect 7 223 17 224
rect 7 211 17 221
rect 428 218 448 225
rect 428 215 448 216
rect 432 211 448 215
rect 7 208 17 209
rect 7 204 13 208
rect 434 195 440 199
rect 430 194 440 195
rect 430 190 440 192
rect 430 186 436 190
rect 48 161 50 165
rect 54 161 58 165
rect 48 159 58 161
rect 48 156 58 157
rect 48 152 54 156
rect 50 144 66 148
rect 46 143 66 144
rect 46 135 66 141
rect 46 132 66 133
rect 46 128 62 132
rect 46 127 66 128
rect 46 118 66 125
rect 46 115 66 116
rect 50 111 66 115
rect 52 95 58 99
rect 48 94 58 95
rect 48 90 58 92
rect 48 86 54 90
rect 8 34 10 38
rect 14 34 18 38
rect 8 33 18 34
rect 8 30 18 31
rect 8 26 14 30
rect 11 9 17 13
rect 7 8 17 9
rect 7 -4 17 6
rect 7 -7 17 -6
rect 7 -11 13 -7
<< pdiffusion >>
rect 9 955 23 959
rect 27 955 29 959
rect 9 953 29 955
rect 9 950 29 951
rect 9 946 25 950
rect 9 945 29 946
rect -7 938 29 942
rect -11 937 29 938
rect 252 936 266 940
rect 270 936 272 940
rect 252 935 272 936
rect -11 934 29 935
rect -11 930 25 934
rect -11 929 29 930
rect 252 932 272 933
rect 256 928 272 932
rect -11 926 29 927
rect -7 922 29 926
rect -11 921 29 922
rect -11 917 29 919
rect -11 913 25 917
rect -11 912 29 913
rect 229 910 265 914
rect -11 909 29 910
rect -7 905 29 909
rect 229 909 269 910
rect 229 905 269 907
rect 233 901 269 905
rect 229 899 269 901
rect 229 896 269 897
rect 9 893 29 894
rect 9 889 25 893
rect 9 888 29 889
rect 229 892 265 896
rect 9 884 29 886
rect 9 880 25 884
rect 233 884 269 888
rect 229 883 269 884
rect 229 879 269 881
rect 233 875 269 879
rect 229 873 269 875
rect 229 869 269 871
rect 229 865 265 869
rect 229 863 269 865
rect 229 859 269 861
rect 233 855 269 859
rect 229 853 269 855
rect 229 850 269 851
rect 229 846 265 850
rect -24 840 -10 844
rect -6 840 -4 844
rect -24 839 -4 840
rect 233 838 269 842
rect -24 836 -4 837
rect -20 832 -4 836
rect 229 837 269 838
rect 229 833 269 835
rect 233 829 269 833
rect 229 827 269 829
rect 229 823 269 825
rect 229 819 265 823
rect -21 815 -5 819
rect -25 814 -5 815
rect 229 817 269 819
rect 391 822 405 826
rect 409 822 411 826
rect 391 820 411 822
rect 391 817 411 818
rect 229 814 269 815
rect -25 809 -5 812
rect -25 805 -10 809
rect -6 805 -5 809
rect -25 802 -5 805
rect 233 810 269 814
rect 391 813 407 817
rect 391 812 411 813
rect 375 805 411 809
rect 371 804 411 805
rect 371 801 411 802
rect -25 799 -5 800
rect -21 795 -5 799
rect 371 797 407 801
rect 371 796 411 797
rect 371 793 411 794
rect 375 789 411 793
rect 371 788 411 789
rect 371 784 411 786
rect 371 780 407 784
rect 371 779 411 780
rect 371 776 411 777
rect 375 772 411 776
rect 9 760 23 764
rect 27 760 29 764
rect 9 758 29 760
rect 391 760 411 761
rect 391 756 407 760
rect 9 755 29 756
rect 9 751 25 755
rect 391 755 411 756
rect 391 751 411 753
rect 9 750 29 751
rect 391 747 407 751
rect -7 743 29 747
rect -11 742 29 743
rect -11 739 29 740
rect -11 735 25 739
rect -11 734 29 735
rect -11 731 29 732
rect -7 727 29 731
rect -11 726 29 727
rect 252 726 266 730
rect 270 726 272 730
rect 252 725 272 726
rect -11 722 29 724
rect -11 718 25 722
rect -11 717 29 718
rect 252 722 272 723
rect 256 718 272 722
rect -11 714 29 715
rect -7 710 29 714
rect 233 700 269 704
rect 9 698 29 699
rect 9 694 25 698
rect 9 693 29 694
rect 229 699 269 700
rect 229 695 269 697
rect 233 691 269 695
rect 9 689 29 691
rect 9 685 25 689
rect 229 689 269 691
rect 229 685 269 687
rect 229 681 265 685
rect 229 679 269 681
rect 229 676 269 677
rect 233 672 269 676
rect 229 664 265 668
rect 229 663 269 664
rect 229 659 269 661
rect 233 655 269 659
rect 229 653 269 655
rect 229 650 269 651
rect 233 646 269 650
rect -24 640 -10 644
rect -6 640 -4 644
rect -24 639 -4 640
rect 229 638 265 642
rect -24 636 -4 637
rect -20 632 -4 636
rect 229 637 269 638
rect 229 633 269 635
rect 233 629 269 633
rect 229 627 269 629
rect 391 628 405 632
rect 409 628 411 632
rect 229 624 269 625
rect 233 620 269 624
rect 391 626 411 628
rect 391 623 411 624
rect 391 619 407 623
rect -21 615 -5 619
rect -25 614 -5 615
rect 391 618 411 619
rect -25 609 -5 612
rect -25 605 -10 609
rect -6 605 -5 609
rect -25 602 -5 605
rect 375 611 411 615
rect 371 610 411 611
rect 371 607 411 608
rect 371 603 407 607
rect -25 599 -5 600
rect -21 595 -5 599
rect 371 602 411 603
rect 371 599 411 600
rect 375 595 411 599
rect 371 594 411 595
rect 371 590 411 592
rect 371 586 407 590
rect 371 585 411 586
rect 371 582 411 583
rect 375 578 411 582
rect 391 566 411 567
rect 9 562 23 566
rect 27 562 29 566
rect 9 560 29 562
rect 391 562 407 566
rect 391 561 411 562
rect 9 557 29 558
rect 9 553 25 557
rect 391 557 411 559
rect 391 553 407 557
rect 9 552 29 553
rect -7 545 29 549
rect -11 544 29 545
rect -11 541 29 542
rect -11 537 25 541
rect -11 536 29 537
rect -11 533 29 534
rect -7 529 29 533
rect -11 528 29 529
rect -11 524 29 526
rect -11 520 25 524
rect -11 519 29 520
rect -11 516 29 517
rect -7 512 29 516
rect 253 505 267 509
rect 271 505 273 509
rect 253 504 273 505
rect 253 501 273 502
rect 9 500 29 501
rect 9 496 25 500
rect 9 495 29 496
rect 257 497 273 501
rect 9 491 29 493
rect 9 487 25 491
rect 236 480 271 485
rect 231 479 271 480
rect 231 476 271 477
rect 235 472 271 476
rect 231 471 271 472
rect 231 468 271 469
rect 231 464 267 468
rect 235 456 271 460
rect 231 455 271 456
rect 231 451 271 453
rect -24 446 -10 450
rect -6 446 -4 450
rect -24 445 -4 446
rect 231 447 267 451
rect -24 442 -4 443
rect -20 438 -4 442
rect 231 445 271 447
rect 231 442 271 443
rect 236 437 271 442
rect 231 435 271 437
rect 231 432 271 433
rect 235 428 271 432
rect -21 421 -5 425
rect -25 420 -5 421
rect -25 415 -5 418
rect -25 411 -10 415
rect -6 411 -5 415
rect -25 408 -5 411
rect 391 415 405 419
rect 409 415 411 419
rect 391 413 411 415
rect 391 410 411 411
rect 391 406 407 410
rect -25 405 -5 406
rect -21 401 -5 405
rect 391 405 411 406
rect 375 398 411 402
rect 371 397 411 398
rect 371 394 411 395
rect 371 390 407 394
rect 371 389 411 390
rect 371 386 411 387
rect 375 382 411 386
rect 371 381 411 382
rect 371 377 411 379
rect 371 373 407 377
rect 371 372 411 373
rect 371 369 411 370
rect 9 364 23 368
rect 27 364 29 368
rect 9 362 29 364
rect 375 365 411 369
rect 9 359 29 360
rect 9 355 25 359
rect 9 354 29 355
rect 391 353 411 354
rect -7 347 29 351
rect -11 346 29 347
rect 391 349 407 353
rect 391 348 411 349
rect 391 344 411 346
rect -11 343 29 344
rect -11 339 25 343
rect -11 338 29 339
rect 391 340 407 344
rect -11 335 29 336
rect -7 331 29 335
rect -11 330 29 331
rect -11 326 29 328
rect -11 322 25 326
rect -11 321 29 322
rect -11 318 29 319
rect -7 314 29 318
rect 9 302 29 303
rect 9 298 25 302
rect 9 297 29 298
rect 253 300 267 304
rect 271 300 273 304
rect 253 299 273 300
rect 253 296 273 297
rect 9 293 29 295
rect 9 289 25 293
rect 257 292 273 296
rect 234 271 270 275
rect 234 270 274 271
rect 234 266 274 268
rect 234 262 270 266
rect 234 260 274 262
rect 391 261 405 265
rect 409 261 411 265
rect 234 256 274 258
rect -24 249 -10 253
rect -6 249 -4 253
rect -24 248 -4 249
rect 238 252 274 256
rect 234 250 274 252
rect 391 259 411 261
rect 391 256 411 257
rect 391 252 407 256
rect 391 251 411 252
rect 234 247 274 248
rect -24 245 -4 246
rect -20 241 -4 245
rect 234 243 270 247
rect 375 244 411 248
rect 371 243 411 244
rect 371 240 411 241
rect 371 236 407 240
rect 371 235 411 236
rect 371 232 411 233
rect 375 228 411 232
rect -21 224 -5 228
rect -25 223 -5 224
rect 371 227 411 228
rect 371 223 411 225
rect -25 218 -5 221
rect -25 214 -10 218
rect -6 214 -5 218
rect -25 211 -5 214
rect 371 219 407 223
rect 371 218 411 219
rect 371 215 411 216
rect 375 211 411 215
rect -25 208 -5 209
rect -21 204 -5 208
rect 391 199 411 200
rect 391 195 407 199
rect 391 194 411 195
rect 391 190 411 192
rect 391 186 407 190
rect 9 161 23 165
rect 27 161 29 165
rect 9 159 29 161
rect 9 156 29 157
rect 9 152 25 156
rect 9 151 29 152
rect -7 144 29 148
rect -11 143 29 144
rect -11 140 29 141
rect -11 136 25 140
rect -11 135 29 136
rect -11 132 29 133
rect -7 128 29 132
rect -11 127 29 128
rect -11 123 29 125
rect -11 119 25 123
rect -11 118 29 119
rect -11 115 29 116
rect -7 111 29 115
rect 9 99 29 100
rect 9 95 25 99
rect 9 94 29 95
rect 9 90 29 92
rect 9 86 25 90
rect -24 34 -10 38
rect -6 34 -4 38
rect -24 33 -4 34
rect -24 30 -4 31
rect -20 26 -4 30
rect -21 9 -5 13
rect -25 8 -5 9
rect -25 3 -5 6
rect -25 -1 -10 3
rect -6 -1 -5 3
rect -25 -4 -5 -1
rect -25 -7 -5 -6
rect -21 -11 -5 -7
<< ndcontact >>
rect 50 955 54 959
rect 54 946 58 950
rect 46 938 50 942
rect 286 936 290 940
rect 290 928 294 932
rect 62 922 66 926
rect 46 905 50 909
rect 283 910 287 914
rect 299 901 303 905
rect 48 889 52 893
rect 299 892 303 896
rect 54 880 58 884
rect 283 884 287 888
rect 299 875 303 879
rect 283 865 287 869
rect 299 855 303 859
rect 299 846 303 850
rect 10 840 14 844
rect 14 832 18 836
rect 283 838 287 842
rect 299 829 303 833
rect 7 815 11 819
rect 432 822 436 826
rect 299 810 303 814
rect 436 813 440 817
rect 428 805 432 809
rect 13 795 17 799
rect 444 789 448 793
rect 428 772 432 776
rect 50 760 54 764
rect 54 751 58 755
rect 430 756 434 760
rect 436 747 440 751
rect 46 743 50 747
rect 62 727 66 731
rect 286 726 290 730
rect 290 718 294 722
rect 46 710 50 714
rect 48 694 52 698
rect 283 700 287 704
rect 54 685 58 689
rect 299 691 303 695
rect 283 672 287 676
rect 283 664 287 668
rect 283 655 287 659
rect 299 646 303 650
rect 10 640 14 644
rect 14 632 18 636
rect 283 638 287 642
rect 283 629 287 633
rect 299 620 303 624
rect 432 628 436 632
rect 436 619 440 623
rect 7 615 11 619
rect 428 611 432 615
rect 13 595 17 599
rect 444 595 448 599
rect 428 578 432 582
rect 50 562 54 566
rect 430 562 434 566
rect 54 553 58 557
rect 436 553 440 557
rect 46 545 50 549
rect 62 529 66 533
rect 46 512 50 516
rect 287 505 291 509
rect 48 496 52 500
rect 291 497 295 501
rect 54 487 58 491
rect 285 480 289 484
rect 301 472 305 476
rect 301 464 305 468
rect 301 456 305 460
rect 10 446 14 450
rect 285 447 289 451
rect 14 438 18 442
rect 285 437 289 441
rect 301 428 305 432
rect 7 421 11 425
rect 432 415 436 419
rect 436 406 440 410
rect 13 401 17 405
rect 428 398 432 402
rect 444 382 448 386
rect 50 364 54 368
rect 428 365 432 369
rect 54 355 58 359
rect 46 347 50 351
rect 430 349 434 353
rect 436 340 440 344
rect 62 331 66 335
rect 46 314 50 318
rect 48 298 52 302
rect 287 300 291 304
rect 54 289 58 293
rect 291 292 295 296
rect 304 271 308 275
rect 288 262 292 266
rect 10 249 14 253
rect 432 261 436 265
rect 436 252 440 256
rect 14 241 18 245
rect 304 243 308 247
rect 428 244 432 248
rect 7 224 11 228
rect 444 228 448 232
rect 428 211 432 215
rect 13 204 17 208
rect 430 195 434 199
rect 436 186 440 190
rect 50 161 54 165
rect 54 152 58 156
rect 46 144 50 148
rect 62 128 66 132
rect 46 111 50 115
rect 48 95 52 99
rect 54 86 58 90
rect 10 34 14 38
rect 14 26 18 30
rect 7 9 11 13
rect 13 -11 17 -7
<< pdcontact >>
rect 23 955 27 959
rect 25 946 29 950
rect -11 938 -7 942
rect 266 936 270 940
rect 25 930 29 934
rect 252 928 256 932
rect -11 922 -7 926
rect 83 922 87 926
rect 25 913 29 917
rect 265 910 269 914
rect -11 905 -7 909
rect 229 901 233 905
rect 25 889 29 893
rect 265 892 269 896
rect 25 880 29 884
rect 229 884 233 888
rect 229 875 233 879
rect 265 865 269 869
rect 229 855 233 859
rect 265 846 269 850
rect -10 840 -6 844
rect 229 838 233 842
rect -24 832 -20 836
rect 229 829 233 833
rect 265 819 269 823
rect -25 815 -21 819
rect 405 822 409 826
rect -10 805 -6 809
rect 229 810 233 814
rect 407 813 411 817
rect 371 805 375 809
rect -25 795 -21 799
rect 407 797 411 801
rect 371 789 375 793
rect 465 789 469 793
rect 407 780 411 784
rect 371 772 375 776
rect 23 760 27 764
rect 407 756 411 760
rect 25 751 29 755
rect 407 747 411 751
rect -11 743 -7 747
rect 25 735 29 739
rect -11 727 -7 731
rect 83 727 87 731
rect 266 726 270 730
rect 25 718 29 722
rect 252 718 256 722
rect -11 710 -7 714
rect 229 700 233 704
rect 25 694 29 698
rect 229 691 233 695
rect 25 685 29 689
rect 265 681 269 685
rect 229 672 233 676
rect 265 664 269 668
rect 229 655 233 659
rect 229 646 233 650
rect -10 640 -6 644
rect 265 638 269 642
rect -24 632 -20 636
rect 229 629 233 633
rect 405 628 409 632
rect 229 620 233 624
rect 407 619 411 623
rect -25 615 -21 619
rect -10 605 -6 609
rect 371 611 375 615
rect 407 603 411 607
rect -25 595 -21 599
rect 371 595 375 599
rect 465 595 469 599
rect 407 586 411 590
rect 371 578 375 582
rect 23 562 27 566
rect 407 562 411 566
rect 25 553 29 557
rect 407 553 411 557
rect -11 545 -7 549
rect 25 537 29 541
rect -11 529 -7 533
rect 83 529 87 533
rect 25 520 29 524
rect -11 512 -7 516
rect 267 505 271 509
rect 25 496 29 500
rect 253 497 257 501
rect 25 487 29 491
rect 231 472 235 476
rect 267 464 271 468
rect 231 456 235 460
rect -10 446 -6 450
rect 267 447 271 451
rect -24 438 -20 442
rect 231 428 235 432
rect -25 421 -21 425
rect -10 411 -6 415
rect 405 415 409 419
rect 407 406 411 410
rect -25 401 -21 405
rect 371 398 375 402
rect 407 390 411 394
rect 371 382 375 386
rect 465 382 469 386
rect 407 373 411 377
rect 23 364 27 368
rect 371 365 375 369
rect 25 355 29 359
rect -11 347 -7 351
rect 407 349 411 353
rect 25 339 29 343
rect 407 340 411 344
rect -11 331 -7 335
rect 83 331 87 335
rect 25 322 29 326
rect -11 314 -7 318
rect 25 298 29 302
rect 267 300 271 304
rect 25 289 29 293
rect 253 292 257 296
rect 270 271 274 275
rect 270 262 274 266
rect 405 261 409 265
rect -10 249 -6 253
rect 234 252 238 256
rect 407 252 411 256
rect -24 241 -20 245
rect 270 243 274 247
rect 371 244 375 248
rect 407 236 411 240
rect 371 228 375 232
rect -25 224 -21 228
rect 465 228 469 232
rect -10 214 -6 218
rect 407 219 411 223
rect 371 211 375 215
rect -25 204 -21 208
rect 407 195 411 199
rect 407 186 411 190
rect 23 161 27 165
rect 25 152 29 156
rect -11 144 -7 148
rect 25 136 29 140
rect -11 128 -7 132
rect 83 128 87 132
rect 25 119 29 123
rect -11 111 -7 115
rect 25 95 29 99
rect 25 86 29 90
rect -10 34 -6 38
rect -24 26 -20 30
rect -25 9 -21 13
rect -10 -1 -6 3
rect -25 -11 -21 -7
<< psubstratepcontact >>
rect 298 928 302 932
rect 70 922 74 926
rect 22 832 26 836
rect 307 810 311 814
rect 21 795 25 799
rect 452 789 456 793
rect 70 727 74 731
rect 298 718 302 722
rect 22 632 26 636
rect 307 628 311 632
rect 21 595 25 599
rect 452 595 456 599
rect 70 529 74 533
rect 299 497 303 501
rect 22 438 26 442
rect 309 432 313 436
rect 21 401 25 405
rect 452 382 456 386
rect 70 331 74 335
rect 299 292 303 296
rect 312 252 316 256
rect 22 241 26 245
rect 452 228 456 232
rect 21 204 25 208
rect 70 128 74 132
rect 22 26 26 30
rect 21 -11 25 -7
<< nsubstratencontact >>
rect 244 928 248 932
rect 25 870 29 874
rect -32 832 -28 836
rect -33 805 -29 809
rect 221 810 225 814
rect 407 737 411 741
rect 244 718 248 722
rect 25 675 29 679
rect -32 632 -28 636
rect 221 620 225 624
rect -33 605 -29 609
rect 407 543 411 547
rect 245 497 249 501
rect 25 477 29 481
rect -32 438 -28 442
rect 223 428 227 432
rect -33 411 -29 415
rect 407 330 411 334
rect 245 292 249 296
rect 25 279 29 283
rect 226 252 230 256
rect -32 241 -28 245
rect -33 214 -29 218
rect 407 176 411 180
rect 25 76 29 80
rect -32 26 -28 30
rect -33 -1 -29 3
<< polysilicon >>
rect 8 951 9 953
rect 29 951 48 953
rect 58 951 61 953
rect -39 935 -11 937
rect 29 935 46 937
rect 66 935 69 937
rect 249 933 252 935
rect 272 933 284 935
rect 294 933 297 935
rect -23 927 -11 929
rect 29 927 46 929
rect 66 927 69 929
rect -40 919 -11 921
rect 29 919 46 921
rect 66 919 69 921
rect -39 910 -11 912
rect 29 910 46 912
rect 66 910 69 912
rect 218 907 229 909
rect 269 907 283 909
rect 303 907 306 909
rect 218 897 229 899
rect 269 897 283 899
rect 303 897 306 899
rect 8 886 9 888
rect 29 886 48 888
rect 58 886 61 888
rect 218 881 229 883
rect 269 881 283 883
rect 303 881 306 883
rect 218 871 229 873
rect 269 871 283 873
rect 303 871 306 873
rect 218 861 229 863
rect 269 861 283 863
rect 303 861 306 863
rect 218 851 229 853
rect 269 851 283 853
rect 303 851 306 853
rect -27 837 -24 839
rect -4 837 8 839
rect 18 837 21 839
rect 218 835 229 837
rect 269 835 283 837
rect 303 835 306 837
rect 218 825 229 827
rect 269 825 283 827
rect 303 825 306 827
rect 390 818 391 820
rect 411 818 430 820
rect 440 818 443 820
rect 218 815 229 817
rect 269 815 283 817
rect 303 815 306 817
rect -36 812 -25 814
rect -5 812 7 814
rect 17 812 20 814
rect -36 800 -25 802
rect -5 800 7 802
rect 17 800 20 802
rect 343 802 371 804
rect 411 802 428 804
rect 448 802 451 804
rect 359 794 371 796
rect 411 794 428 796
rect 448 794 451 796
rect 342 786 371 788
rect 411 786 428 788
rect 448 786 451 788
rect 343 777 371 779
rect 411 777 428 779
rect 448 777 451 779
rect 8 756 9 758
rect 29 756 48 758
rect 58 756 61 758
rect 390 753 391 755
rect 411 753 430 755
rect 440 753 443 755
rect -39 740 -11 742
rect 29 740 46 742
rect 66 740 69 742
rect -23 732 -11 734
rect 29 732 46 734
rect 66 732 69 734
rect -40 724 -11 726
rect 29 724 46 726
rect 66 724 69 726
rect 249 723 252 725
rect 272 723 284 725
rect 294 723 297 725
rect -39 715 -11 717
rect 29 715 46 717
rect 66 715 69 717
rect 218 697 229 699
rect 269 697 283 699
rect 303 697 306 699
rect 8 691 9 693
rect 29 691 48 693
rect 58 691 61 693
rect 218 687 229 689
rect 269 687 283 689
rect 303 687 306 689
rect 218 677 229 679
rect 269 677 283 679
rect 303 677 306 679
rect 218 661 229 663
rect 269 661 283 663
rect 303 661 306 663
rect 218 651 229 653
rect 269 651 283 653
rect 303 651 306 653
rect -27 637 -24 639
rect -4 637 8 639
rect 18 637 21 639
rect 218 635 229 637
rect 269 635 283 637
rect 303 635 306 637
rect 218 625 229 627
rect 269 625 283 627
rect 303 625 306 627
rect 390 624 391 626
rect 411 624 430 626
rect 440 624 443 626
rect -36 612 -25 614
rect -5 612 7 614
rect 17 612 20 614
rect 343 608 371 610
rect 411 608 428 610
rect 448 608 451 610
rect -36 600 -25 602
rect -5 600 7 602
rect 17 600 20 602
rect 359 600 371 602
rect 411 600 428 602
rect 448 600 451 602
rect 342 592 371 594
rect 411 592 428 594
rect 448 592 451 594
rect 343 583 371 585
rect 411 583 428 585
rect 448 583 451 585
rect 8 558 9 560
rect 29 558 48 560
rect 58 558 61 560
rect 390 559 391 561
rect 411 559 430 561
rect 440 559 443 561
rect -39 542 -11 544
rect 29 542 46 544
rect 66 542 69 544
rect -23 534 -11 536
rect 29 534 46 536
rect 66 534 69 536
rect -40 526 -11 528
rect 29 526 46 528
rect 66 526 69 528
rect -39 517 -11 519
rect 29 517 46 519
rect 66 517 69 519
rect 250 502 253 504
rect 273 502 285 504
rect 295 502 298 504
rect 8 493 9 495
rect 29 493 48 495
rect 58 493 61 495
rect 219 477 231 479
rect 271 477 285 479
rect 305 477 308 479
rect 219 469 231 471
rect 271 469 285 471
rect 305 469 308 471
rect 219 453 231 455
rect 271 453 285 455
rect 305 453 308 455
rect -27 443 -24 445
rect -4 443 8 445
rect 18 443 21 445
rect 219 443 231 445
rect 271 443 285 445
rect 305 443 308 445
rect 219 433 231 435
rect 271 433 285 435
rect 305 433 308 435
rect -36 418 -25 420
rect -5 418 7 420
rect 17 418 20 420
rect 390 411 391 413
rect 411 411 430 413
rect 440 411 443 413
rect -36 406 -25 408
rect -5 406 7 408
rect 17 406 20 408
rect 343 395 371 397
rect 411 395 428 397
rect 448 395 451 397
rect 359 387 371 389
rect 411 387 428 389
rect 448 387 451 389
rect 342 379 371 381
rect 411 379 428 381
rect 448 379 451 381
rect 343 370 371 372
rect 411 370 428 372
rect 448 370 451 372
rect 8 360 9 362
rect 29 360 48 362
rect 58 360 61 362
rect -39 344 -11 346
rect 29 344 46 346
rect 66 344 69 346
rect 390 346 391 348
rect 411 346 430 348
rect 440 346 443 348
rect -23 336 -11 338
rect 29 336 46 338
rect 66 336 69 338
rect -40 328 -11 330
rect 29 328 46 330
rect 66 328 69 330
rect -39 319 -11 321
rect 29 319 46 321
rect 66 319 69 321
rect 250 297 253 299
rect 273 297 285 299
rect 295 297 298 299
rect 8 295 9 297
rect 29 295 48 297
rect 58 295 61 297
rect 223 268 234 270
rect 274 268 288 270
rect 308 268 311 270
rect 223 258 234 260
rect 274 258 288 260
rect 308 258 311 260
rect -27 246 -24 248
rect -4 246 8 248
rect 18 246 21 248
rect 390 257 391 259
rect 411 257 430 259
rect 440 257 443 259
rect 223 248 234 250
rect 274 248 288 250
rect 308 248 311 250
rect 343 241 371 243
rect 411 241 428 243
rect 448 241 451 243
rect 359 233 371 235
rect 411 233 428 235
rect 448 233 451 235
rect 342 225 371 227
rect 411 225 428 227
rect 448 225 451 227
rect -36 221 -25 223
rect -5 221 7 223
rect 17 221 20 223
rect 343 216 371 218
rect 411 216 428 218
rect 448 216 451 218
rect -36 209 -25 211
rect -5 209 7 211
rect 17 209 20 211
rect 390 192 391 194
rect 411 192 430 194
rect 440 192 443 194
rect 8 157 9 159
rect 29 157 48 159
rect 58 157 61 159
rect -39 141 -11 143
rect 29 141 46 143
rect 66 141 69 143
rect -23 133 -11 135
rect 29 133 46 135
rect 66 133 69 135
rect -40 125 -11 127
rect 29 125 46 127
rect 66 125 69 127
rect -39 116 -11 118
rect 29 116 46 118
rect 66 116 69 118
rect 8 92 9 94
rect 29 92 48 94
rect 58 92 61 94
rect -27 31 -24 33
rect -4 31 8 33
rect 18 31 21 33
rect -36 6 -25 8
rect -5 6 7 8
rect 17 6 20 8
rect -36 -6 -25 -4
rect -5 -6 7 -4
rect 17 -6 20 -4
<< polycontact >>
rect 4 950 8 954
rect -43 934 -39 938
rect -27 926 -23 930
rect 275 929 279 933
rect -44 918 -40 922
rect -43 909 -39 913
rect 214 906 218 910
rect 214 896 218 900
rect 4 885 8 889
rect 214 880 218 884
rect 214 870 218 874
rect 214 860 218 864
rect 214 850 218 854
rect -1 833 3 837
rect 214 834 218 838
rect 214 824 218 828
rect -40 811 -36 815
rect 214 814 218 818
rect 386 817 390 821
rect -40 799 -36 803
rect 339 801 343 805
rect 355 793 359 797
rect 338 785 342 789
rect 339 776 343 780
rect 4 755 8 759
rect 386 752 390 756
rect -43 739 -39 743
rect -27 731 -23 735
rect -44 723 -40 727
rect -43 714 -39 718
rect 275 719 279 723
rect 4 690 8 694
rect 214 696 218 700
rect 214 686 218 690
rect 214 676 218 680
rect 214 660 218 664
rect 214 650 218 654
rect -1 633 3 637
rect 214 634 218 638
rect 214 624 218 628
rect 386 623 390 627
rect -40 611 -36 615
rect -40 599 -36 603
rect 339 607 343 611
rect 355 599 359 603
rect 338 591 342 595
rect 339 582 343 586
rect 4 557 8 561
rect 386 558 390 562
rect -43 541 -39 545
rect -27 533 -23 537
rect -44 525 -40 529
rect -43 516 -39 520
rect 4 492 8 496
rect 276 498 280 502
rect 215 476 219 480
rect 215 468 219 472
rect 215 452 219 456
rect -1 439 3 443
rect 215 442 219 446
rect 215 432 219 436
rect -40 417 -36 421
rect -40 405 -36 409
rect 386 410 390 414
rect 339 394 343 398
rect 355 386 359 390
rect 338 378 342 382
rect 339 369 343 373
rect 4 359 8 363
rect -43 343 -39 347
rect 386 345 390 349
rect -27 335 -23 339
rect -44 327 -40 331
rect -43 318 -39 322
rect 4 294 8 298
rect 276 293 280 297
rect 219 267 223 271
rect 219 257 223 261
rect 219 247 223 251
rect 386 256 390 260
rect -1 242 3 246
rect 339 240 343 244
rect 355 232 359 236
rect -40 220 -36 224
rect 338 224 342 228
rect -40 208 -36 212
rect 339 215 343 219
rect 386 191 390 195
rect 4 156 8 160
rect -43 140 -39 144
rect -27 132 -23 136
rect -44 124 -40 128
rect -43 115 -39 119
rect 4 91 8 95
rect -1 27 3 31
rect -40 5 -36 9
rect -40 -7 -36 -3
<< metal1 >>
rect -43 962 36 966
rect -43 938 -39 962
rect 32 959 36 962
rect 27 955 50 959
rect -35 950 4 954
rect -44 922 -40 925
rect -35 913 -31 950
rect 29 946 32 950
rect 58 946 74 950
rect -19 938 -11 942
rect -39 909 -31 913
rect -27 901 -23 926
rect -19 926 -15 938
rect 41 934 45 938
rect 29 930 45 934
rect -19 922 -11 926
rect -19 909 -15 922
rect 29 913 32 917
rect 41 909 45 930
rect 70 926 74 946
rect 66 922 70 926
rect 74 922 83 926
rect -19 905 -11 909
rect 41 905 46 909
rect -27 897 44 901
rect 40 893 44 897
rect 29 889 48 893
rect -31 885 4 889
rect 29 880 32 884
rect 70 884 74 922
rect 58 880 74 884
rect 25 874 29 880
rect -1 844 3 847
rect -6 840 10 844
rect -28 832 -24 836
rect -1 819 3 833
rect 18 832 22 836
rect -33 815 -25 819
rect -1 815 7 819
rect -44 811 -40 815
rect -33 809 -29 815
rect -1 809 3 815
rect -6 805 3 809
rect -44 799 -40 803
rect -33 799 -29 805
rect -33 795 -25 799
rect 17 795 21 799
rect -43 767 36 771
rect -43 743 -39 767
rect 32 764 36 767
rect 27 760 50 764
rect -35 755 4 759
rect -44 727 -40 730
rect -35 718 -31 755
rect 29 751 32 755
rect 58 751 74 755
rect -19 743 -11 747
rect -39 714 -31 718
rect -27 706 -23 731
rect -19 731 -15 743
rect 41 739 45 743
rect 29 735 45 739
rect -19 727 -11 731
rect -19 714 -15 727
rect 29 718 32 722
rect 41 714 45 735
rect 70 731 74 751
rect 66 727 70 731
rect 74 727 83 731
rect -19 710 -11 714
rect 41 710 46 714
rect -27 702 44 706
rect 40 698 44 702
rect 29 694 48 698
rect -31 690 4 694
rect 29 685 32 689
rect 70 689 74 727
rect 58 685 74 689
rect 25 679 29 685
rect -1 644 3 647
rect -6 640 10 644
rect -28 632 -24 636
rect -1 619 3 633
rect 18 632 22 636
rect -33 615 -25 619
rect -1 615 7 619
rect -44 611 -40 615
rect -33 609 -29 615
rect -1 609 3 615
rect -6 605 3 609
rect -44 599 -40 603
rect -33 599 -29 605
rect -33 595 -25 599
rect 17 595 21 599
rect -43 569 36 573
rect -43 545 -39 569
rect 32 566 36 569
rect 27 562 50 566
rect -35 557 4 561
rect -44 529 -40 532
rect -35 520 -31 557
rect 29 553 32 557
rect 58 553 74 557
rect -19 545 -11 549
rect -39 516 -31 520
rect -27 508 -23 533
rect -19 533 -15 545
rect 41 541 45 545
rect 29 537 45 541
rect -19 529 -11 533
rect -19 516 -15 529
rect 29 520 32 524
rect 41 516 45 537
rect 70 533 74 553
rect 66 529 70 533
rect 74 529 83 533
rect -19 512 -11 516
rect 41 512 46 516
rect -27 504 44 508
rect 40 500 44 504
rect 29 496 48 500
rect -31 492 4 496
rect 29 487 32 491
rect 70 491 74 529
rect 58 487 74 491
rect 25 481 29 487
rect -1 450 3 453
rect -6 446 10 450
rect -28 438 -24 442
rect -1 425 3 439
rect 18 438 22 442
rect -33 421 -25 425
rect -1 421 7 425
rect -44 417 -40 421
rect -33 415 -29 421
rect -1 415 3 421
rect -6 411 3 415
rect -44 405 -40 409
rect -33 405 -29 411
rect -33 401 -25 405
rect 17 401 21 405
rect -43 371 36 375
rect -43 347 -39 371
rect 32 368 36 371
rect 27 364 50 368
rect -35 359 4 363
rect -44 331 -40 334
rect -35 322 -31 359
rect 29 355 32 359
rect 58 355 74 359
rect -19 347 -11 351
rect -39 318 -31 322
rect -27 310 -23 335
rect -19 335 -15 347
rect 41 343 45 347
rect 29 339 45 343
rect -19 331 -11 335
rect -19 318 -15 331
rect 29 322 32 326
rect 41 318 45 339
rect 70 335 74 355
rect 66 331 70 335
rect 74 331 83 335
rect -19 314 -11 318
rect 41 314 46 318
rect -27 306 44 310
rect 40 302 44 306
rect 29 298 48 302
rect -31 294 4 298
rect 29 289 32 293
rect 70 293 74 331
rect 58 289 74 293
rect 25 283 29 289
rect -1 253 3 256
rect -6 249 10 253
rect -28 241 -24 245
rect -1 228 3 242
rect 18 241 22 245
rect -33 224 -25 228
rect -1 224 7 228
rect -44 220 -40 224
rect -33 218 -29 224
rect -1 218 3 224
rect -6 214 3 218
rect -44 208 -40 212
rect -33 208 -29 214
rect -33 204 -25 208
rect 17 204 21 208
rect -43 168 36 172
rect -43 144 -39 168
rect 32 165 36 168
rect 27 161 50 165
rect -35 156 4 160
rect -44 128 -40 131
rect -35 119 -31 156
rect 29 152 32 156
rect 58 152 74 156
rect -19 144 -11 148
rect -39 115 -31 119
rect -27 107 -23 132
rect -19 132 -15 144
rect 41 140 45 144
rect 29 136 45 140
rect -19 128 -11 132
rect -19 115 -15 128
rect 29 119 32 123
rect 41 115 45 136
rect 70 132 74 152
rect 66 128 70 132
rect 74 128 83 132
rect -19 111 -11 115
rect 41 111 46 115
rect -27 103 44 107
rect 40 99 44 103
rect 29 95 48 99
rect -31 91 4 95
rect 29 86 32 90
rect 70 90 74 128
rect 58 86 74 90
rect 25 80 29 86
rect -1 38 3 41
rect -6 34 10 38
rect -28 26 -24 30
rect -1 13 3 27
rect 18 26 22 30
rect -33 9 -25 13
rect -1 9 7 13
rect -44 5 -40 9
rect -33 3 -29 9
rect -1 3 3 9
rect -6 -1 3 3
rect -44 -7 -40 -3
rect -33 -7 -29 -1
rect -33 -11 -25 -7
rect 17 -11 21 -7
rect 107 -32 111 993
rect 115 819 119 993
rect 123 855 127 993
rect 115 691 119 814
rect 123 701 127 850
rect 131 829 135 993
rect 139 865 143 993
rect 115 472 119 686
rect 123 481 127 696
rect 131 681 135 824
rect 115 252 119 467
rect 123 272 127 476
rect 131 457 135 676
rect 139 655 143 860
rect 147 839 151 993
rect 155 901 159 993
rect 147 665 151 834
rect 131 375 135 452
rect 139 437 143 650
rect 147 577 151 660
rect 155 629 159 896
rect 163 875 167 993
rect 171 911 175 993
rect 179 970 183 993
rect 179 885 183 965
rect 163 775 167 870
rect 179 797 183 880
rect 163 639 167 770
rect 163 603 167 634
rect 147 447 151 572
rect 147 390 151 442
rect 131 262 135 370
rect 115 220 119 247
rect 131 236 135 257
rect 115 46 119 215
rect 187 -32 191 993
rect 275 940 279 943
rect 270 936 286 940
rect 248 928 252 932
rect 275 914 279 929
rect 294 928 298 932
rect 269 910 283 914
rect 212 906 214 910
rect 212 896 214 900
rect 229 888 233 901
rect 212 880 214 884
rect 221 875 229 879
rect 212 870 214 874
rect 212 860 214 864
rect 212 850 214 854
rect 212 834 214 838
rect 221 833 225 875
rect 265 869 269 892
rect 277 888 281 910
rect 303 901 311 905
rect 277 884 283 888
rect 299 879 303 892
rect 229 842 233 855
rect 221 829 229 833
rect 212 824 214 828
rect 212 814 214 818
rect 221 814 225 829
rect 265 823 269 846
rect 283 842 287 865
rect 307 859 311 901
rect 303 855 311 859
rect 299 833 303 846
rect 307 814 311 855
rect 225 810 229 814
rect 303 810 307 814
rect 339 829 418 833
rect 339 805 343 829
rect 414 826 418 829
rect 409 822 432 826
rect 347 817 386 821
rect 338 789 342 792
rect 347 780 351 817
rect 411 813 414 817
rect 440 813 456 817
rect 363 805 371 809
rect 338 776 339 780
rect 343 776 351 780
rect 355 768 359 793
rect 363 793 367 805
rect 423 801 427 805
rect 411 797 427 801
rect 363 789 371 793
rect 363 776 367 789
rect 411 780 414 784
rect 423 776 427 797
rect 452 793 456 813
rect 448 789 452 793
rect 456 789 465 793
rect 363 772 371 776
rect 423 772 428 776
rect 355 764 426 768
rect 422 760 426 764
rect 411 756 430 760
rect 351 752 386 756
rect 411 747 414 751
rect 452 751 456 789
rect 440 747 456 751
rect 407 741 411 747
rect 275 730 279 733
rect 270 726 286 730
rect 248 718 252 722
rect 221 700 229 704
rect 212 696 214 700
rect 212 686 214 690
rect 212 676 214 680
rect 212 660 214 664
rect 221 659 225 700
rect 229 676 233 691
rect 275 685 279 719
rect 294 718 298 722
rect 269 681 279 685
rect 275 668 279 681
rect 269 664 279 668
rect 283 676 287 700
rect 303 691 311 695
rect 283 668 287 672
rect 221 655 229 659
rect 212 650 214 654
rect 212 634 214 638
rect 229 633 233 646
rect 275 642 279 664
rect 269 638 279 642
rect 283 642 287 655
rect 307 650 311 691
rect 303 646 311 650
rect 275 633 279 638
rect 275 629 283 633
rect 307 632 311 646
rect 212 624 214 628
rect 307 624 311 628
rect 225 620 229 624
rect 303 620 311 624
rect 339 635 418 639
rect 339 611 343 635
rect 414 632 418 635
rect 409 628 432 632
rect 347 623 386 627
rect 338 595 342 598
rect 347 586 351 623
rect 411 619 414 623
rect 440 619 456 623
rect 363 611 371 615
rect 338 582 339 586
rect 343 582 351 586
rect 355 574 359 599
rect 363 599 367 611
rect 423 607 427 611
rect 411 603 427 607
rect 363 595 371 599
rect 363 582 367 595
rect 411 586 414 590
rect 423 582 427 603
rect 452 599 456 619
rect 448 595 452 599
rect 456 595 465 599
rect 363 578 371 582
rect 423 578 428 582
rect 355 570 426 574
rect 422 566 426 570
rect 411 562 430 566
rect 351 558 386 562
rect 411 553 414 557
rect 452 557 456 595
rect 440 553 456 557
rect 407 547 411 553
rect 276 509 280 512
rect 271 505 287 509
rect 249 497 253 501
rect 212 476 215 480
rect 212 468 215 472
rect 231 460 235 472
rect 276 468 280 498
rect 295 497 299 501
rect 271 464 280 468
rect 212 452 215 456
rect 276 451 280 464
rect 271 447 280 451
rect 285 451 289 480
rect 305 472 313 476
rect 301 460 305 464
rect 212 442 215 446
rect 276 441 280 447
rect 276 437 285 441
rect 309 436 313 472
rect 212 432 215 436
rect 227 428 231 432
rect 305 428 313 432
rect 339 422 418 426
rect 339 398 343 422
rect 414 419 418 422
rect 409 415 432 419
rect 347 410 386 414
rect 338 382 342 385
rect 347 373 351 410
rect 411 406 414 410
rect 440 406 456 410
rect 363 398 371 402
rect 338 369 339 373
rect 343 369 351 373
rect 355 361 359 386
rect 363 386 367 398
rect 423 394 427 398
rect 411 390 427 394
rect 363 382 371 386
rect 363 369 367 382
rect 411 373 414 377
rect 423 369 427 390
rect 452 386 456 406
rect 448 382 452 386
rect 456 382 465 386
rect 363 365 371 369
rect 423 365 428 369
rect 355 357 426 361
rect 422 353 426 357
rect 411 349 430 353
rect 351 345 386 349
rect 411 340 414 344
rect 452 344 456 382
rect 440 340 456 344
rect 407 334 411 340
rect 276 304 280 307
rect 271 300 287 304
rect 249 292 253 296
rect 276 275 280 293
rect 295 292 299 296
rect 274 271 287 275
rect 308 271 316 275
rect 212 267 219 271
rect 283 266 287 271
rect 274 262 279 266
rect 283 262 288 266
rect 212 257 219 261
rect 230 252 234 256
rect 212 247 219 251
rect 275 247 279 262
rect 312 256 316 271
rect 312 247 316 252
rect 274 243 279 247
rect 308 243 316 247
rect 339 268 418 272
rect 339 244 343 268
rect 414 265 418 268
rect 409 261 432 265
rect 347 256 386 260
rect 338 228 342 231
rect 347 219 351 256
rect 411 252 414 256
rect 440 252 456 256
rect 363 244 371 248
rect 338 215 339 219
rect 343 215 351 219
rect 355 207 359 232
rect 363 232 367 244
rect 423 240 427 244
rect 411 236 427 240
rect 363 228 371 232
rect 363 215 367 228
rect 411 219 414 223
rect 423 215 427 236
rect 452 232 456 252
rect 448 228 452 232
rect 456 228 465 232
rect 363 211 371 215
rect 423 211 428 215
rect 355 203 426 207
rect 422 199 426 203
rect 411 195 430 199
rect 351 191 386 195
rect 411 186 414 190
rect 452 190 456 228
rect 440 186 456 190
rect 407 180 411 186
<< m2contact >>
rect -45 925 -40 930
rect 32 945 37 950
rect 41 938 46 943
rect 32 913 37 918
rect -36 885 -31 890
rect 32 880 37 885
rect -1 847 4 852
rect -45 730 -40 735
rect 32 750 37 755
rect 41 743 46 748
rect 32 718 37 723
rect -36 690 -31 695
rect 32 685 37 690
rect -1 647 4 652
rect -45 532 -40 537
rect 32 552 37 557
rect 41 545 46 550
rect 32 520 37 525
rect -36 492 -31 497
rect 32 487 37 492
rect -1 453 4 458
rect -45 334 -40 339
rect 32 354 37 359
rect 41 347 46 352
rect 32 322 37 327
rect -36 294 -31 299
rect 32 289 37 294
rect -1 256 4 261
rect -45 131 -40 136
rect 32 151 37 156
rect 41 144 46 149
rect 32 119 37 124
rect -36 91 -31 96
rect 32 86 37 91
rect -1 41 4 46
rect 123 850 128 855
rect 115 814 120 819
rect 139 860 144 865
rect 131 824 136 829
rect 123 696 128 701
rect 115 686 120 691
rect 131 676 136 681
rect 123 476 128 481
rect 115 467 120 472
rect 155 896 160 901
rect 147 834 152 839
rect 147 660 152 665
rect 139 650 144 655
rect 131 452 136 457
rect 178 965 183 970
rect 171 906 176 911
rect 179 880 184 885
rect 163 870 168 875
rect 179 792 184 797
rect 162 770 167 775
rect 163 634 168 639
rect 155 624 160 629
rect 163 598 168 603
rect 146 572 151 577
rect 147 442 152 447
rect 139 432 144 437
rect 147 385 152 390
rect 130 370 135 375
rect 123 267 128 272
rect 131 257 136 262
rect 115 247 120 252
rect 131 231 136 236
rect 115 215 120 220
rect 114 41 119 46
rect 275 943 280 948
rect 207 906 212 911
rect 207 896 212 901
rect 207 880 212 885
rect 207 870 212 875
rect 207 860 212 865
rect 207 850 212 855
rect 207 834 212 839
rect 207 824 212 829
rect 207 814 212 819
rect 337 792 342 797
rect 333 776 338 781
rect 414 812 419 817
rect 423 805 428 810
rect 414 780 419 785
rect 346 752 351 757
rect 414 747 419 752
rect 275 733 280 738
rect 207 696 212 701
rect 207 686 212 691
rect 207 676 212 681
rect 207 660 212 665
rect 207 650 212 655
rect 207 634 212 639
rect 207 624 212 629
rect 337 598 342 603
rect 333 582 338 587
rect 414 618 419 623
rect 423 611 428 616
rect 414 586 419 591
rect 346 558 351 563
rect 414 553 419 558
rect 276 512 281 517
rect 207 476 212 481
rect 207 467 212 472
rect 207 452 212 457
rect 207 442 212 447
rect 207 432 212 437
rect 337 385 342 390
rect 333 369 338 374
rect 414 405 419 410
rect 423 398 428 403
rect 414 373 419 378
rect 346 345 351 350
rect 414 340 419 345
rect 276 307 281 312
rect 207 267 212 272
rect 207 257 212 262
rect 207 247 212 252
rect 337 231 342 236
rect 333 215 338 220
rect 414 251 419 256
rect 423 244 428 249
rect 414 219 419 224
rect 346 191 351 196
rect 414 186 419 191
<< pdm12contact >>
rect 231 480 236 485
rect 231 437 236 442
<< metal2 >>
rect 41 965 178 970
rect -40 926 -31 930
rect -36 890 -31 926
rect 33 918 37 945
rect 41 943 46 965
rect 280 943 322 948
rect 33 885 37 913
rect 96 906 171 911
rect 176 906 207 911
rect 96 852 101 906
rect 160 896 207 901
rect 184 880 207 885
rect 168 870 207 875
rect 144 860 207 865
rect 4 847 101 852
rect 128 850 207 855
rect 152 834 207 839
rect 423 835 460 840
rect 136 824 207 829
rect 120 814 207 819
rect 184 792 337 797
rect 342 793 351 797
rect 275 776 333 781
rect 41 770 162 775
rect -40 731 -31 735
rect -36 695 -31 731
rect 33 723 37 750
rect 41 748 46 770
rect 275 738 280 776
rect 346 757 351 793
rect 415 785 419 812
rect 423 810 428 835
rect 415 752 419 780
rect 33 690 37 718
rect 128 696 207 701
rect 120 686 207 691
rect 136 676 207 681
rect 152 660 207 665
rect 4 647 50 652
rect 144 650 207 655
rect 45 629 50 647
rect 423 641 460 646
rect 168 634 207 639
rect 45 624 155 629
rect 160 624 207 629
rect 168 598 337 603
rect 342 599 351 603
rect 276 582 333 587
rect 41 572 146 577
rect -40 533 -31 537
rect -36 497 -31 533
rect 33 525 37 552
rect 41 550 46 572
rect 33 492 37 520
rect 276 517 281 582
rect 346 563 351 599
rect 415 591 419 618
rect 423 616 428 641
rect 415 558 419 586
rect 128 476 207 481
rect 224 480 231 485
rect 120 467 207 472
rect 4 453 70 458
rect 65 437 70 453
rect 136 452 207 457
rect 152 442 207 447
rect 224 442 229 480
rect 224 437 231 442
rect 65 432 139 437
rect 144 432 207 437
rect 423 428 460 433
rect 152 385 337 390
rect 342 386 351 390
rect 41 370 130 375
rect -40 335 -31 339
rect -36 299 -31 335
rect 33 327 37 354
rect 41 352 46 370
rect 276 369 333 374
rect 33 294 37 322
rect 276 312 281 369
rect 346 350 351 386
rect 415 378 419 405
rect 423 403 428 428
rect 415 345 419 373
rect 423 274 460 279
rect -1 267 123 272
rect 128 267 207 272
rect -1 261 4 267
rect 136 257 207 262
rect 120 247 207 252
rect 136 231 337 236
rect 342 232 351 236
rect 120 215 333 220
rect 346 196 351 232
rect 415 224 419 251
rect 423 249 428 274
rect 415 191 419 219
rect 41 166 345 171
rect -40 132 -31 136
rect -36 96 -31 132
rect 33 124 37 151
rect 41 149 46 166
rect 33 91 37 119
rect 4 41 114 46
<< labels >>
rlabel metal1 116 992 118 993 5 G0
rlabel metal1 124 992 126 993 5 G1
rlabel metal1 132 992 134 993 5 P1
rlabel metal1 140 992 142 993 5 G2
rlabel metal1 148 992 150 993 5 P2
rlabel metal1 156 992 158 993 5 G3
rlabel metal1 164 992 166 993 5 P3
rlabel metal1 172 992 174 993 5 G4
rlabel metal1 180 992 182 993 5 P4
rlabel metal1 276 921 278 922 7 C5_bar
rlabel metal1 297 928 298 932 7 gnd
rlabel metal1 249 928 250 932 7 vdd
rlabel polycontact 214 907 215 909 7 G4
rlabel polycontact 214 897 215 899 7 G3
rlabel polycontact 214 881 215 883 7 P4
rlabel polycontact 214 871 215 873 7 P3
rlabel polycontact 214 861 215 863 7 G2
rlabel polycontact 214 851 215 853 7 G1
rlabel polycontact 214 835 215 837 7 P2
rlabel polycontact 214 825 215 827 7 P1
rlabel polycontact 214 815 215 817 7 G0
rlabel psubstratepcontact 307 810 311 814 7 gnd
rlabel nsubstratencontact 222 811 223 813 7 vdd
rlabel metal1 276 711 278 712 7 C4_bar
rlabel metal1 297 718 298 722 7 gnd
rlabel metal1 249 718 250 722 7 vdd
rlabel polycontact 214 697 215 699 3 G1
rlabel polycontact 214 687 215 689 3 G0
rlabel polycontact 214 677 215 679 3 P1
rlabel polycontact 214 661 215 663 3 P2
rlabel polycontact 214 651 215 653 3 G2
rlabel polycontact 214 635 215 637 3 P3
rlabel polycontact 214 625 215 627 3 G3
rlabel nsubstratencontact 222 621 224 623 7 vdd
rlabel metal1 308 620 310 623 8 gnd
rlabel metal1 277 490 279 491 7 C3_bar
rlabel metal1 298 497 299 501 7 gnd
rlabel metal1 250 497 251 501 7 vdd
rlabel metal1 213 477 214 479 3 G1
rlabel metal1 213 469 214 471 3 G0
rlabel metal1 213 453 214 455 3 P1
rlabel metal1 213 443 214 445 3 P2
rlabel metal1 213 433 214 435 3 G2
rlabel nsubstratencontact 226 429 227 431 7 vdd
rlabel metal1 310 428 311 430 7 gnd
rlabel metal1 226 252 227 255 3 vdd
rlabel metal1 217 247 218 250 3 G0
rlabel metal1 217 267 218 270 3 G1
rlabel metal1 250 292 251 296 7 vdd
rlabel metal1 298 292 299 296 7 gnd
rlabel metal1 278 279 279 284 7 C2_bar
rlabel metal1 313 243 314 246 8 gnd
rlabel metal1 217 257 218 260 3 P1
rlabel polycontact -44 918 -40 922 1 B4
rlabel polycontact -43 909 -39 913 1 A4
rlabel metal1 61 946 62 950 7 gnd
rlabel nsubstratencontact 25 870 29 874 1 vdd
rlabel metal1 1 822 2 827 1 G4_bar
rlabel metal1 -44 812 -43 814 1 B4
rlabel metal1 -44 800 -43 802 1 A4
rlabel metal1 21 832 22 836 7 gnd
rlabel metal1 -27 832 -26 836 7 vdd
rlabel metal1 -33 795 -32 799 3 vdd
rlabel metal1 19 795 21 796 8 gnd
rlabel polycontact -44 723 -40 727 1 B3
rlabel polycontact -43 714 -39 718 1 A3
rlabel metal1 68 727 74 731 7 gnd
rlabel metal1 61 751 62 755 7 gnd
rlabel nsubstratencontact 25 675 29 679 1 vdd
rlabel metal1 1 622 2 627 1 G3_bar
rlabel metal1 -44 612 -43 614 1 B3
rlabel metal1 -44 600 -43 602 1 A3
rlabel metal1 21 632 22 636 7 gnd
rlabel metal1 -27 632 -26 636 7 vdd
rlabel metal1 -33 595 -32 599 3 vdd
rlabel metal1 19 595 21 596 8 gnd
rlabel nsubstratencontact 25 477 29 481 1 vdd
rlabel metal1 61 553 62 557 7 gnd
rlabel metal1 68 529 74 533 7 gnd
rlabel polycontact -43 516 -39 520 3 A2
rlabel polycontact -44 525 -40 529 3 B2
rlabel metal1 19 401 21 402 8 gnd
rlabel metal1 -33 401 -32 405 3 vdd
rlabel metal1 -27 438 -26 442 7 vdd
rlabel metal1 21 438 22 442 7 gnd
rlabel metal1 -44 406 -43 408 1 A2
rlabel metal1 -44 418 -43 420 1 B2
rlabel metal1 1 428 2 433 1 G2_bar
rlabel polycontact -44 327 -40 331 3 B1
rlabel polycontact -43 318 -39 322 3 A1
rlabel nsubstratencontact 25 279 29 283 1 vdd
rlabel metal1 61 355 62 359 7 gnd
rlabel metal1 68 331 74 335 7 gnd
rlabel metal1 1 231 2 236 1 G1_bar
rlabel metal1 -44 221 -43 223 3 A1
rlabel metal1 -44 209 -43 211 3 B1
rlabel metal1 21 241 22 245 7 gnd
rlabel metal1 -27 241 -26 245 7 vdd
rlabel metal1 -33 204 -32 208 3 vdd
rlabel metal1 19 204 21 205 8 gnd
rlabel polycontact -44 124 -40 128 3 B0
rlabel polycontact -43 115 -39 119 3 A0
rlabel nsubstratencontact 25 76 29 80 1 vdd
rlabel metal1 61 152 62 156 7 gnd
rlabel metal1 68 128 74 132 7 gnd
rlabel metal1 21 26 22 30 7 gnd
rlabel metal1 -27 26 -26 30 7 vdd
rlabel metal1 -33 -11 -32 -7 3 vdd
rlabel metal1 19 -11 21 -10 8 gnd
rlabel metal1 -44 -6 -43 -4 1 A0
rlabel metal1 -44 6 -43 8 1 B0
rlabel metal1 1 16 2 21 1 G0_bar
rlabel polycontact 338 224 342 228 1 P1
rlabel metal1 450 228 456 232 7 gnd
rlabel metal1 443 252 444 256 7 gnd
rlabel nsubstratencontact 407 176 411 180 1 vdd
rlabel nsubstratencontact 407 330 411 334 1 vdd
rlabel metal1 443 406 444 410 7 gnd
rlabel metal1 450 382 456 386 7 gnd
rlabel metal1 450 595 456 599 7 gnd
rlabel metal1 443 619 444 623 7 gnd
rlabel nsubstratencontact 407 543 411 547 1 vdd
rlabel nsubstratencontact 407 737 411 741 1 vdd
rlabel metal1 443 813 444 817 7 gnd
rlabel metal1 450 789 456 793 7 gnd
rlabel polycontact 339 215 343 219 1 G0
rlabel polycontact 339 369 343 373 1 C2
rlabel polycontact 338 378 342 382 1 P2
rlabel polycontact 339 582 343 586 1 C3
rlabel polycontact 338 591 342 595 1 P3
rlabel polycontact 339 776 343 780 1 C4
rlabel polycontact 338 785 342 789 1 P4
rlabel metal2 426 837 429 839 1 S4
rlabel metal2 426 642 429 644 1 S3
rlabel metal2 425 429 428 431 1 S2
rlabel metal2 426 276 429 278 1 S1
rlabel metal2 333 168 336 170 1 S0
rlabel metal2 313 944 321 946 1 C5
<< end >>
